LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

-- Top Block --
ENTITY c_10bit2char_vga_H256 IS --chinese
PORT(
	X0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X4 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X5 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X6 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X7 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X8 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X9 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X10 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X11 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X12 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X13 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X14 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X15 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	
	Y0 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	Y1 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	Y2 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	Y3 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	Y4 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	Y5 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	Y6 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	Y7 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	Y8 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	Y9 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	Y10 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	Y11 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	Y12 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	Y13 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	Y14 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	Y15 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000");	
END c_10bit2char_vga_H256;

ARCHITECTURE convert OF c_10bit2char_vga_H256 IS
	BEGIN
		Y0 <= X0;
		Y1 <= X1;
		Y2 <= X2;
		Y3 <= X3;
		Y4 <= X4;
		Y5 <= X5;
		Y6 <= X6;
		Y7 <= X7;
		Y8 <= X8;
		Y9 <= X9;
		Y10 <= X10;
		Y11 <= X11;
		Y12 <= X12;
		Y13 <= X13;
		Y14 <= X14;
		Y15 <= X15;
END convert;