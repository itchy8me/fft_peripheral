-- *************************************************************************
-- Author : Wernher Korff																	*
-- Function : follows clock signal when ready is '1' and converting is '0'	*
-- *************************************************************************

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY convert2spectrum IS
	PORT(
		-- R is real and I is imaginary
		X0R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X0I: IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X3R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X3I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X4R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X4I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X5R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X5I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X6R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X6I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X7R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X7I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X8R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X8I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X9R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X9I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X10R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X10I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X11R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X11I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X12R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X12I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X13R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X13I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X14R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X14I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X15R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X15I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		
		incoming128set : IN STD_LOGIC := '0';
		
		converting : OUT STD_LOGIC := '0');
END clock_control;