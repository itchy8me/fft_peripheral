-- *************************************************************************
-- Author : Wernher Korff																	*
-- Function : shift 2048 samples into fft												*
-- *************************************************************************

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
--USE IEEE.STD_LOGIC_ARITH.ALL;


--Shifts in 8 samples for parallel data ouput N=8 big
ENTITY c_2048to16x128_shifter IS
	PORT(
			--X0 downto X2048 ports input from ADC	
		X0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X4 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X5 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X6 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X7 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X8 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X9 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X10 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X11 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X12 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X13 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X14 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X15 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X16 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X17 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X18 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X19 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X20 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X21 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X22 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X23 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X24 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X25 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X26 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X27 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X28 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X29 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X30 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X31 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X32 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X33 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X34 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X35 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X36 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X37 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X38 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X39 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X40 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X41 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X42 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X43 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X44 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X45 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X46 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X47 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X48 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X49 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X50 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X51 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X52 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X53 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X54 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X55 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X56 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X57 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X58 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X59 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X60 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X61 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X62 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X63 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X64 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X65 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X66 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X67 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X68 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X69 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X70 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X71 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X72 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X73 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X74 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X75 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X76 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X77 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X78 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X79 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X80 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X81 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X82 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X83 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X84 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X85 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X86 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X87 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X88 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X89 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X90 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X91 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X92 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X93 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X94 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X95 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X96 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X97 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X98 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X99 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X100 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X101 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X102 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X103 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X104 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X105 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X106 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X107 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X108 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X109 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X110 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X111 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X112 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X113 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X114 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X115 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X116 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X117 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X118 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X119 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X120 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X121 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X122 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X123 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X124 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X125 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X126 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X127 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X128 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X129 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X130 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X131 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X132 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X133 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X134 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X135 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X136 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X137 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X138 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X139 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X140 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X141 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X142 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X143 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X144 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X145 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X146 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X147 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X148 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X149 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X150 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X151 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X152 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X153 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X154 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X155 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X156 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X157 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X158 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X159 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X160 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X161 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X162 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X163 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X164 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X165 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X166 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X167 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X168 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X169 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X170 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X171 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X172 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X173 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X174 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X175 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X176 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X177 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X178 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X179 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X180 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X181 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X182 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X183 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X184 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X185 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X186 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X187 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X188 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X189 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X190 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X191 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X192 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X193 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X194 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X195 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X196 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X197 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X198 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X199 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X200 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X201 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X202 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X203 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X204 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X205 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X206 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X207 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X208 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X209 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X210 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X211 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X212 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X213 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X214 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X215 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X216 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X217 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X218 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X219 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X220 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X221 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X222 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X223 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X224 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X225 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X226 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X227 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X228 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X229 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X230 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X231 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X232 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X233 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X234 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X235 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X236 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X237 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X238 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X239 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X240 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X241 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X242 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X243 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X244 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X245 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X246 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X247 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X248 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X249 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X250 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X251 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X252 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X253 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X254 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X255 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X256 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X257 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X258 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X259 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X260 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X261 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X262 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X263 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X264 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X265 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X266 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X267 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X268 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X269 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X270 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X271 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X272 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X273 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X274 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X275 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X276 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X277 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X278 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X279 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X280 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X281 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X282 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X283 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X284 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X285 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X286 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X287 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X288 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X289 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X290 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X291 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X292 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X293 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X294 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X295 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X296 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X297 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X298 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X299 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X300 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X301 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X302 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X303 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X304 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X305 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X306 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X307 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X308 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X309 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X310 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X311 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X312 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X313 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X314 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X315 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X316 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X317 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X318 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X319 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X320 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X321 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X322 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X323 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X324 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X325 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X326 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X327 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X328 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X329 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X330 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X331 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X332 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X333 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X334 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X335 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X336 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X337 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X338 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X339 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X340 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X341 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X342 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X343 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X344 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X345 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X346 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X347 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X348 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X349 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X350 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X351 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X352 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X353 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X354 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X355 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X356 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X357 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X358 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X359 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X360 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X361 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X362 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X363 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X364 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X365 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X366 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X367 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X368 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X369 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X370 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X371 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X372 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X373 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X374 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X375 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X376 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X377 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X378 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X379 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X380 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X381 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X382 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X383 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X384 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X385 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X386 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X387 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X388 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X389 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X390 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X391 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X392 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X393 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X394 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X395 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X396 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X397 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X398 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X399 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X400 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X401 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X402 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X403 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X404 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X405 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X406 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X407 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X408 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X409 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X410 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X411 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X412 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X413 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X414 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X415 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X416 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X417 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X418 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X419 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X420 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X421 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X422 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X423 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X424 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X425 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X426 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X427 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X428 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X429 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X430 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X431 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X432 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X433 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X434 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X435 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X436 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X437 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X438 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X439 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X440 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X441 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X442 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X443 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X444 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X445 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X446 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X447 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X448 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X449 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X450 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X451 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X452 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X453 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X454 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X455 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X456 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X457 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X458 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X459 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X460 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X461 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X462 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X463 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X464 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X465 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X466 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X467 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X468 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X469 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X470 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X471 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X472 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X473 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X474 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X475 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X476 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X477 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X478 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X479 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X480 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X481 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X482 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X483 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X484 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X485 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X486 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X487 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X488 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X489 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X490 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X491 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X492 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X493 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X494 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X495 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X496 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X497 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X498 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X499 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X500 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X501 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X502 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X503 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X504 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X505 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X506 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X507 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X508 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X509 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X510 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X511 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X512 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X513 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X514 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X515 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X516 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X517 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X518 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X519 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X520 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X521 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X522 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X523 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X524 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X525 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X526 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X527 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X528 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X529 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X530 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X531 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X532 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X533 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X534 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X535 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X536 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X537 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X538 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X539 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X540 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X541 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X542 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X543 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X544 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X545 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X546 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X547 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X548 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X549 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X550 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X551 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X552 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X553 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X554 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X555 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X556 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X557 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X558 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X559 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X560 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X561 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X562 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X563 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X564 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X565 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X566 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X567 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X568 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X569 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X570 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X571 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X572 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X573 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X574 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X575 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X576 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X577 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X578 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X579 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X580 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X581 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X582 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X583 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X584 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X585 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X586 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X587 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X588 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X589 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X590 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X591 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X592 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X593 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X594 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X595 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X596 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X597 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X598 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X599 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X600 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X601 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X602 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X603 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X604 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X605 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X606 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X607 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X608 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X609 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X610 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X611 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X612 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X613 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X614 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X615 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X616 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X617 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X618 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X619 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X620 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X621 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X622 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X623 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X624 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X625 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X626 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X627 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X628 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X629 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X630 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X631 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X632 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X633 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X634 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X635 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X636 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X637 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X638 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X639 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X640 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X641 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X642 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X643 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X644 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X645 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X646 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X647 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X648 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X649 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X650 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X651 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X652 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X653 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X654 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X655 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X656 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X657 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X658 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X659 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X660 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X661 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X662 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X663 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X664 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X665 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X666 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X667 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X668 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X669 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X670 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X671 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X672 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X673 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X674 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X675 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X676 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X677 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X678 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X679 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X680 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X681 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X682 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X683 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X684 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X685 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X686 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X687 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X688 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X689 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X690 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X691 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X692 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X693 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X694 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X695 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X696 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X697 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X698 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X699 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X700 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X701 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X702 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X703 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X704 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X705 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X706 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X707 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X708 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X709 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X710 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X711 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X712 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X713 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X714 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X715 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X716 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X717 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X718 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X719 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X720 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X721 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X722 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X723 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X724 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X725 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X726 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X727 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X728 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X729 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X730 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X731 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X732 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X733 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X734 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X735 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X736 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X737 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X738 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X739 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X740 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X741 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X742 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X743 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X744 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X745 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X746 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X747 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X748 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X749 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X750 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X751 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X752 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X753 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X754 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X755 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X756 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X757 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X758 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X759 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X760 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X761 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X762 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X763 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X764 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X765 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X766 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X767 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X768 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X769 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X770 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X771 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X772 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X773 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X774 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X775 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X776 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X777 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X778 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X779 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X780 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X781 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X782 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X783 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X784 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X785 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X786 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X787 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X788 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X789 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X790 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X791 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X792 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X793 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X794 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X795 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X796 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X797 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X798 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X799 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X800 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X801 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X802 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X803 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X804 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X805 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X806 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X807 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X808 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X809 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X810 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X811 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X812 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X813 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X814 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X815 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X816 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X817 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X818 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X819 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X820 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X821 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X822 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X823 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X824 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X825 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X826 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X827 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X828 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X829 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X830 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X831 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X832 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X833 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X834 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X835 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X836 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X837 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X838 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X839 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X840 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X841 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X842 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X843 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X844 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X845 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X846 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X847 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X848 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X849 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X850 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X851 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X852 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X853 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X854 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X855 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X856 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X857 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X858 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X859 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X860 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X861 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X862 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X863 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X864 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X865 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X866 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X867 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X868 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X869 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X870 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X871 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X872 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X873 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X874 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X875 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X876 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X877 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X878 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X879 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X880 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X881 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X882 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X883 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X884 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X885 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X886 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X887 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X888 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X889 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X890 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X891 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X892 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X893 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X894 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X895 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X896 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X897 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X898 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X899 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X900 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X901 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X902 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X903 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X904 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X905 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X906 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X907 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X908 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X909 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X910 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X911 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X912 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X913 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X914 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X915 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X916 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X917 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X918 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X919 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X920 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X921 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X922 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X923 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X924 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X925 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X926 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X927 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X928 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X929 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X930 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X931 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X932 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X933 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X934 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X935 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X936 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X937 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X938 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X939 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X940 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X941 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X942 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X943 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X944 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X945 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X946 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X947 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X948 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X949 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X950 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X951 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X952 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X953 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X954 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X955 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X956 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X957 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X958 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X959 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X960 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X961 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X962 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X963 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X964 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X965 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X966 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X967 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X968 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X969 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X970 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X971 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X972 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X973 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X974 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X975 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X976 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X977 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X978 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X979 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X980 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X981 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X982 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X983 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X984 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X985 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X986 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X987 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X988 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X989 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X990 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X991 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X992 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X993 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X994 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X995 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X996 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X997 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X998 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X999 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1000 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1001 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1002 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1003 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1004 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1005 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1006 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1007 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1008 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1009 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1010 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1011 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1012 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1013 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1014 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1015 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1016 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1017 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1018 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1019 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1020 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1021 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1022 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1023 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1024 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1025 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1026 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1027 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1028 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1029 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1030 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1031 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1032 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1033 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1034 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1035 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1036 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1037 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1038 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1039 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1040 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1041 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1042 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1043 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1044 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1045 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1046 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1047 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1048 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1049 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1050 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1051 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1052 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1053 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1054 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1055 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1056 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1057 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1058 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1059 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1060 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1061 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1062 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1063 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1064 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1065 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1066 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1067 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1068 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1069 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1070 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1071 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1072 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1073 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1074 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1075 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1076 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1077 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1078 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1079 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1080 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1081 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1082 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1083 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1084 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1085 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1086 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1087 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1088 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1089 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1090 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1091 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1092 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1093 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1094 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1095 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1096 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1097 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1098 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1099 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1100 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1101 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1102 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1103 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1104 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1105 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1106 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1107 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1108 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1109 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1110 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1111 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1112 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1113 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1114 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1115 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1116 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1117 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1118 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1119 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1120 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1121 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1122 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1123 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1124 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1125 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1126 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1127 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1128 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1129 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1130 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1131 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1132 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1133 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1134 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1135 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1136 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1137 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1138 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1139 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1140 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1141 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1142 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1143 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1144 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1145 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1146 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1147 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1148 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1149 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1150 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1151 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1152 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1153 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1154 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1155 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1156 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1157 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1158 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1159 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1160 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1161 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1162 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1163 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1164 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1165 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1166 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1167 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1168 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1169 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1170 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1171 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1172 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1173 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1174 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1175 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1176 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1177 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1178 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1179 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1180 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1181 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1182 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1183 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1184 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1185 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1186 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1187 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1188 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1189 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1190 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1191 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1192 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1193 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1194 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1195 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1196 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1197 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1198 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1199 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1200 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1201 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1202 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1203 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1204 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1205 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1206 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1207 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1208 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1209 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1210 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1211 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1212 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1213 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1214 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1215 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1216 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1217 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1218 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1219 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1220 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1221 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1222 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1223 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1224 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1225 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1226 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1227 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1228 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1229 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1230 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1231 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1232 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1233 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1234 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1235 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1236 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1237 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1238 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1239 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1240 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1241 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1242 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1243 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1244 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1245 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1246 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1247 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1248 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1249 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1250 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1251 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1252 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1253 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1254 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1255 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1256 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1257 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1258 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1259 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1260 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1261 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1262 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1263 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1264 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1265 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1266 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1267 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1268 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1269 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1270 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1271 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1272 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1273 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1274 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1275 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1276 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1277 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1278 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1279 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1280 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1281 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1282 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1283 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1284 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1285 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1286 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1287 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1288 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1289 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1290 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1291 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1292 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1293 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1294 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1295 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1296 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1297 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1298 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1299 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1300 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1301 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1302 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1303 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1304 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1305 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1306 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1307 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1308 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1309 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1310 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1311 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1312 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1313 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1314 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1315 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1316 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1317 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1318 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1319 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1320 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1321 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1322 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1323 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1324 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1325 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1326 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1327 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1328 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1329 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1330 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1331 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1332 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1333 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1334 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1335 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1336 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1337 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1338 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1339 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1340 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1341 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1342 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1343 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1344 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1345 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1346 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1347 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1348 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1349 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1350 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1351 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1352 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1353 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1354 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1355 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1356 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1357 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1358 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1359 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1360 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1361 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1362 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1363 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1364 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1365 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1366 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1367 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1368 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1369 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1370 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1371 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1372 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1373 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1374 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1375 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1376 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1377 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1378 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1379 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1380 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1381 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1382 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1383 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1384 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1385 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1386 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1387 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1388 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1389 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1390 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1391 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1392 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1393 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1394 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1395 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1396 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1397 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1398 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1399 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1400 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1401 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1402 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1403 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1404 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1405 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1406 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1407 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1408 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1409 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1410 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1411 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1412 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1413 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1414 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1415 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1416 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1417 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1418 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1419 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1420 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1421 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1422 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1423 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1424 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1425 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1426 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1427 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1428 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1429 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1430 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1431 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1432 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1433 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1434 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1435 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1436 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1437 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1438 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1439 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1440 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1441 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1442 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1443 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1444 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1445 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1446 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1447 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1448 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1449 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1450 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1451 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1452 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1453 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1454 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1455 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1456 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1457 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1458 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1459 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1460 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1461 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1462 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1463 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1464 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1465 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1466 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1467 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1468 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1469 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1470 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1471 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1472 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1473 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1474 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1475 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1476 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1477 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1478 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1479 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1480 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1481 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1482 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1483 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1484 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1485 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1486 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1487 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1488 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1489 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1490 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1491 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1492 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1493 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1494 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1495 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1496 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1497 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1498 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1499 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1500 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1501 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1502 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1503 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1504 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1505 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1506 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1507 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1508 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1509 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1510 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1511 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1512 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1513 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1514 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1515 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1516 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1517 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1518 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1519 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1520 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1521 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1522 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1523 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1524 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1525 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1526 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1527 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1528 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1529 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1530 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1531 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1532 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1533 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1534 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1535 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1536 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1537 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1538 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1539 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1540 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1541 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1542 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1543 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1544 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1545 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1546 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1547 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1548 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1549 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1550 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1551 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1552 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1553 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1554 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1555 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1556 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1557 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1558 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1559 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1560 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1561 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1562 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1563 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1564 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1565 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1566 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1567 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1568 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1569 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1570 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1571 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1572 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1573 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1574 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1575 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1576 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1577 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1578 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1579 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1580 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1581 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1582 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1583 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1584 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1585 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1586 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1587 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1588 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1589 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1590 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1591 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1592 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1593 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1594 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1595 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1596 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1597 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1598 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1599 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1600 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1601 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1602 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1603 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1604 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1605 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1606 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1607 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1608 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1609 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1610 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1611 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1612 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1613 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1614 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1615 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1616 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1617 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1618 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1619 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1620 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1621 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1622 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1623 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1624 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1625 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1626 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1627 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1628 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1629 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1630 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1631 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1632 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1633 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1634 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1635 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1636 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1637 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1638 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1639 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1640 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1641 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1642 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1643 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1644 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1645 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1646 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1647 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1648 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1649 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1650 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1651 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1652 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1653 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1654 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1655 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1656 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1657 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1658 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1659 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1660 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1661 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1662 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1663 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1664 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1665 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1666 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1667 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1668 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1669 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1670 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1671 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1672 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1673 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1674 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1675 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1676 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1677 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1678 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1679 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1680 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1681 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1682 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1683 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1684 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1685 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1686 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1687 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1688 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1689 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1690 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1691 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1692 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1693 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1694 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1695 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1696 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1697 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1698 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1699 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1700 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1701 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1702 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1703 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1704 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1705 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1706 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1707 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1708 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1709 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1710 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1711 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1712 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1713 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1714 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1715 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1716 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1717 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1718 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1719 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1720 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1721 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1722 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1723 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1724 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1725 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1726 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1727 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1728 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1729 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1730 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1731 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1732 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1733 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1734 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1735 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1736 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1737 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1738 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1739 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1740 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1741 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1742 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1743 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1744 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1745 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1746 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1747 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1748 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1749 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1750 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1751 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1752 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1753 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1754 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1755 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1756 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1757 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1758 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1759 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1760 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1761 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1762 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1763 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1764 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1765 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1766 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1767 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1768 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1769 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1770 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1771 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1772 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1773 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1774 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1775 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1776 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1777 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1778 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1779 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1780 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1781 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1782 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1783 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1784 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1785 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1786 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1787 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1788 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1789 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1790 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1791 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1792 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1793 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1794 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1795 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1796 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1797 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1798 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1799 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1800 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1801 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1802 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1803 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1804 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1805 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1806 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1807 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1808 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1809 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1810 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1811 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1812 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1813 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1814 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1815 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1816 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1817 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1818 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1819 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1820 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1821 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1822 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1823 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1824 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1825 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1826 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1827 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1828 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1829 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1830 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1831 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1832 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1833 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1834 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1835 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1836 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1837 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1838 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1839 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1840 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1841 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1842 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1843 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1844 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1845 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1846 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1847 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1848 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1849 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1850 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1851 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1852 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1853 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1854 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1855 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1856 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1857 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1858 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1859 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1860 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1861 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1862 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1863 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1864 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1865 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1866 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1867 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1868 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1869 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1870 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1871 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1872 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1873 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1874 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1875 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1876 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1877 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1878 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1879 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1880 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1881 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1882 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1883 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1884 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1885 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1886 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1887 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1888 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1889 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1890 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1891 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1892 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1893 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1894 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1895 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1896 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1897 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1898 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1899 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1900 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1901 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1902 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1903 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1904 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1905 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1906 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1907 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1908 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1909 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1910 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1911 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1912 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1913 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1914 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1915 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1916 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1917 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1918 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1919 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1920 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1921 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1922 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1923 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1924 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1925 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1926 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1927 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1928 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1929 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1930 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1931 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1932 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1933 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1934 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1935 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1936 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1937 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1938 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1939 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1940 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1941 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1942 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1943 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1944 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1945 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1946 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1947 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1948 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1949 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1950 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1951 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1952 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1953 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1954 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1955 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1956 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1957 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1958 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1959 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1960 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1961 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1962 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1963 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1964 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1965 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1966 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1967 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1968 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1969 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1970 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1971 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1972 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1973 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1974 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1975 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1976 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1977 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1978 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1979 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1980 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1981 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1982 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1983 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1984 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1985 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1986 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1987 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1988 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1989 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1990 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1991 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1992 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1993 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1994 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1995 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1996 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1997 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1998 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1999 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2000 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2001 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2002 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2003 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2004 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2005 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2006 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2007 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2008 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2009 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2010 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2011 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2012 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2013 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2014 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2015 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2016 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2017 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2018 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2019 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2020 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2021 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2022 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2023 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2024 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2025 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2026 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2027 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2028 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2029 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2030 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2031 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2032 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2033 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2034 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2035 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2036 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2037 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2038 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2039 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2040 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2041 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2042 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2043 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2044 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2045 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2046 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2047 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		
		-- enable : IN STD_LOGIC := '0';
		fft_finished : IN STD_LOGIC := '0';
		samples_ready : IN STD_LOGIC := '0';
		clk : IN STD_LOGIC := '0';
		
		-- sig_next : OUT STD_LOGIC := '0';
		shift_out0 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out1 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out2 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out3 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out4 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out5 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out6 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out7 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out8 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out9 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out10 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out11 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out12 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out13 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out14 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out15 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000");
END c_2048to16x128_shifter;


--the 4 bit to 7 bit (hex representation) decoding
ARCHITECTURE shift OF c_2048to16x128_shifter IS
	SIGNAL i : INTEGER := 0;
	SIGNAL reading_input : INTEGER := 0;
	-- SIGNAL data_incoming : STD_LOGIC := '0';
		
	BEGIN

	PROCESS(clk,samples_ready,reading_input)
		BEGIN
			
			IF rising_edge(clk) THEN
			IF (samples_ready = '1') THEN
				reading_input <= 1;
			END IF;
			
			IF (fft_finished = '1') THEN
			END IF;
			
			CASE reading_input IS	-- shift the 2048 samples into the FFT
			WHEN 1 =>
					ASE i IS
					WHEN 0 =>
						shift_out0 <= X0;
						shift_out1 <= X1;
						shift_out2 <= X2;
						shift_out3 <= X3;
						shift_out4 <= X4;
						shift_out5 <= X5;
						shift_out6 <= X6;
						shift_out7 <= X7;
						shift_out8 <= X8;
						shift_out9 <= X9;
						shift_out10 <= X10;
						shift_out11 <= X11;
						shift_out12 <= X12;
						shift_out13 <= X13;
						shift_out14 <= X14;
						shift_out15 <= X15;
						i <= i + 1;
					WHEN 1 =>
						shift_out0 <= X16;
						shift_out1 <= X17;
						shift_out2 <= X18;
						shift_out3 <= X19;
						shift_out4 <= X20;
						shift_out5 <= X21;
						shift_out6 <= X22;
						shift_out7 <= X23;
						shift_out8 <= X24;
						shift_out9 <= X25;
						shift_out10 <= X26;
						shift_out11 <= X27;
						shift_out12 <= X28;
						shift_out13 <= X29;
						shift_out14 <= X30;
						shift_out15 <= X31;
						i <= i + 1;
					WHEN 2 =>
						shift_out0 <= X32;
						shift_out1 <= X33;
						shift_out2 <= X34;
						shift_out3 <= X35;
						shift_out4 <= X36;
						shift_out5 <= X37;
						shift_out6 <= X38;
						shift_out7 <= X39;
						shift_out8 <= X40;
						shift_out9 <= X41;
						shift_out10 <= X42;
						shift_out11 <= X43;
						shift_out12 <= X44;
						shift_out13 <= X45;
						shift_out14 <= X46;
						shift_out15 <= X47;
						i <= i + 1;
					WHEN 3 =>
						shift_out0 <= X48;
						shift_out1 <= X49;
						shift_out2 <= X50;
						shift_out3 <= X51;
						shift_out4 <= X52;
						shift_out5 <= X53;
						shift_out6 <= X54;
						shift_out7 <= X55;
						shift_out8 <= X56;
						shift_out9 <= X57;
						shift_out10 <= X58;
						shift_out11 <= X59;
						shift_out12 <= X60;
						shift_out13 <= X61;
						shift_out14 <= X62;
						shift_out15 <= X63;
						i <= i + 1;
					WHEN 4 =>
						shift_out0 <= X64;
						shift_out1 <= X65;
						shift_out2 <= X66;
						shift_out3 <= X67;
						shift_out4 <= X68;
						shift_out5 <= X69;
						shift_out6 <= X70;
						shift_out7 <= X71;
						shift_out8 <= X72;
						shift_out9 <= X73;
						shift_out10 <= X74;
						shift_out11 <= X75;
						shift_out12 <= X76;
						shift_out13 <= X77;
						shift_out14 <= X78;
						shift_out15 <= X79;
						i <= i + 1;
					WHEN 5 =>
						shift_out0 <= X80;
						shift_out1 <= X81;
						shift_out2 <= X82;
						shift_out3 <= X83;
						shift_out4 <= X84;
						shift_out5 <= X85;
						shift_out6 <= X86;
						shift_out7 <= X87;
						shift_out8 <= X88;
						shift_out9 <= X89;
						shift_out10 <= X90;
						shift_out11 <= X91;
						shift_out12 <= X92;
						shift_out13 <= X93;
						shift_out14 <= X94;
						shift_out15 <= X95;
						i <= i + 1;
					WHEN 6 =>
						shift_out0 <= X96;
						shift_out1 <= X97;
						shift_out2 <= X98;
						shift_out3 <= X99;
						shift_out4 <= X100;
						shift_out5 <= X101;
						shift_out6 <= X102;
						shift_out7 <= X103;
						shift_out8 <= X104;
						shift_out9 <= X105;
						shift_out10 <= X106;
						shift_out11 <= X107;
						shift_out12 <= X108;
						shift_out13 <= X109;
						shift_out14 <= X110;
						shift_out15 <= X111;
						i <= i + 1;
					WHEN 7 =>
						shift_out0 <= X112;
						shift_out1 <= X113;
						shift_out2 <= X114;
						shift_out3 <= X115;
						shift_out4 <= X116;
						shift_out5 <= X117;
						shift_out6 <= X118;
						shift_out7 <= X119;
						shift_out8 <= X120;
						shift_out9 <= X121;
						shift_out10 <= X122;
						shift_out11 <= X123;
						shift_out12 <= X124;
						shift_out13 <= X125;
						shift_out14 <= X126;
						shift_out15 <= X127;
						i <= i + 1;
					WHEN 8 =>
						shift_out0 <= X128;
						shift_out1 <= X129;
						shift_out2 <= X130;
						shift_out3 <= X131;
						shift_out4 <= X132;
						shift_out5 <= X133;
						shift_out6 <= X134;
						shift_out7 <= X135;
						shift_out8 <= X136;
						shift_out9 <= X137;
						shift_out10 <= X138;
						shift_out11 <= X139;
						shift_out12 <= X140;
						shift_out13 <= X141;
						shift_out14 <= X142;
						shift_out15 <= X143;
						i <= i + 1;
					WHEN 9 =>
						shift_out0 <= X144;
						shift_out1 <= X145;
						shift_out2 <= X146;
						shift_out3 <= X147;
						shift_out4 <= X148;
						shift_out5 <= X149;
						shift_out6 <= X150;
						shift_out7 <= X151;
						shift_out8 <= X152;
						shift_out9 <= X153;
						shift_out10 <= X154;
						shift_out11 <= X155;
						shift_out12 <= X156;
						shift_out13 <= X157;
						shift_out14 <= X158;
						shift_out15 <= X159;
						i <= i + 1;
					WHEN 10 =>
						shift_out0 <= X160;
						shift_out1 <= X161;
						shift_out2 <= X162;
						shift_out3 <= X163;
						shift_out4 <= X164;
						shift_out5 <= X165;
						shift_out6 <= X166;
						shift_out7 <= X167;
						shift_out8 <= X168;
						shift_out9 <= X169;
						shift_out10 <= X170;
						shift_out11 <= X171;
						shift_out12 <= X172;
						shift_out13 <= X173;
						shift_out14 <= X174;
						shift_out15 <= X175;
						i <= i + 1;
					WHEN 11 =>
						shift_out0 <= X176;
						shift_out1 <= X177;
						shift_out2 <= X178;
						shift_out3 <= X179;
						shift_out4 <= X180;
						shift_out5 <= X181;
						shift_out6 <= X182;
						shift_out7 <= X183;
						shift_out8 <= X184;
						shift_out9 <= X185;
						shift_out10 <= X186;
						shift_out11 <= X187;
						shift_out12 <= X188;
						shift_out13 <= X189;
						shift_out14 <= X190;
						shift_out15 <= X191;
						i <= i + 1;
					WHEN 12 =>
						shift_out0 <= X192;
						shift_out1 <= X193;
						shift_out2 <= X194;
						shift_out3 <= X195;
						shift_out4 <= X196;
						shift_out5 <= X197;
						shift_out6 <= X198;
						shift_out7 <= X199;
						shift_out8 <= X200;
						shift_out9 <= X201;
						shift_out10 <= X202;
						shift_out11 <= X203;
						shift_out12 <= X204;
						shift_out13 <= X205;
						shift_out14 <= X206;
						shift_out15 <= X207;
						i <= i + 1;
					WHEN 13 =>
						shift_out0 <= X208;
						shift_out1 <= X209;
						shift_out2 <= X210;
						shift_out3 <= X211;
						shift_out4 <= X212;
						shift_out5 <= X213;
						shift_out6 <= X214;
						shift_out7 <= X215;
						shift_out8 <= X216;
						shift_out9 <= X217;
						shift_out10 <= X218;
						shift_out11 <= X219;
						shift_out12 <= X220;
						shift_out13 <= X221;
						shift_out14 <= X222;
						shift_out15 <= X223;
						i <= i + 1;
					WHEN 14 =>
						shift_out0 <= X224;
						shift_out1 <= X225;
						shift_out2 <= X226;
						shift_out3 <= X227;
						shift_out4 <= X228;
						shift_out5 <= X229;
						shift_out6 <= X230;
						shift_out7 <= X231;
						shift_out8 <= X232;
						shift_out9 <= X233;
						shift_out10 <= X234;
						shift_out11 <= X235;
						shift_out12 <= X236;
						shift_out13 <= X237;
						shift_out14 <= X238;
						shift_out15 <= X239;
						i <= i + 1;
					WHEN 15 =>
						shift_out0 <= X240;
						shift_out1 <= X241;
						shift_out2 <= X242;
						shift_out3 <= X243;
						shift_out4 <= X244;
						shift_out5 <= X245;
						shift_out6 <= X246;
						shift_out7 <= X247;
						shift_out8 <= X248;
						shift_out9 <= X249;
						shift_out10 <= X250;
						shift_out11 <= X251;
						shift_out12 <= X252;
						shift_out13 <= X253;
						shift_out14 <= X254;
						shift_out15 <= X255;
						i <= i + 1;
					WHEN 16 =>
						shift_out0 <= X256;
						shift_out1 <= X257;
						shift_out2 <= X258;
						shift_out3 <= X259;
						shift_out4 <= X260;
						shift_out5 <= X261;
						shift_out6 <= X262;
						shift_out7 <= X263;
						shift_out8 <= X264;
						shift_out9 <= X265;
						shift_out10 <= X266;
						shift_out11 <= X267;
						shift_out12 <= X268;
						shift_out13 <= X269;
						shift_out14 <= X270;
						shift_out15 <= X271;
						i <= i + 1;
					WHEN 17 =>
						shift_out0 <= X272;
						shift_out1 <= X273;
						shift_out2 <= X274;
						shift_out3 <= X275;
						shift_out4 <= X276;
						shift_out5 <= X277;
						shift_out6 <= X278;
						shift_out7 <= X279;
						shift_out8 <= X280;
						shift_out9 <= X281;
						shift_out10 <= X282;
						shift_out11 <= X283;
						shift_out12 <= X284;
						shift_out13 <= X285;
						shift_out14 <= X286;
						shift_out15 <= X287;
						i <= i + 1;
					WHEN 18 =>
						shift_out0 <= X288;
						shift_out1 <= X289;
						shift_out2 <= X290;
						shift_out3 <= X291;
						shift_out4 <= X292;
						shift_out5 <= X293;
						shift_out6 <= X294;
						shift_out7 <= X295;
						shift_out8 <= X296;
						shift_out9 <= X297;
						shift_out10 <= X298;
						shift_out11 <= X299;
						shift_out12 <= X300;
						shift_out13 <= X301;
						shift_out14 <= X302;
						shift_out15 <= X303;
						i <= i + 1;
					WHEN 19 =>
						shift_out0 <= X304;
						shift_out1 <= X305;
						shift_out2 <= X306;
						shift_out3 <= X307;
						shift_out4 <= X308;
						shift_out5 <= X309;
						shift_out6 <= X310;
						shift_out7 <= X311;
						shift_out8 <= X312;
						shift_out9 <= X313;
						shift_out10 <= X314;
						shift_out11 <= X315;
						shift_out12 <= X316;
						shift_out13 <= X317;
						shift_out14 <= X318;
						shift_out15 <= X319;
						i <= i + 1;
					WHEN 20 =>
						shift_out0 <= X320;
						shift_out1 <= X321;
						shift_out2 <= X322;
						shift_out3 <= X323;
						shift_out4 <= X324;
						shift_out5 <= X325;
						shift_out6 <= X326;
						shift_out7 <= X327;
						shift_out8 <= X328;
						shift_out9 <= X329;
						shift_out10 <= X330;
						shift_out11 <= X331;
						shift_out12 <= X332;
						shift_out13 <= X333;
						shift_out14 <= X334;
						shift_out15 <= X335;
						i <= i + 1;
					WHEN 21 =>
						shift_out0 <= X336;
						shift_out1 <= X337;
						shift_out2 <= X338;
						shift_out3 <= X339;
						shift_out4 <= X340;
						shift_out5 <= X341;
						shift_out6 <= X342;
						shift_out7 <= X343;
						shift_out8 <= X344;
						shift_out9 <= X345;
						shift_out10 <= X346;
						shift_out11 <= X347;
						shift_out12 <= X348;
						shift_out13 <= X349;
						shift_out14 <= X350;
						shift_out15 <= X351;
						i <= i + 1;
					WHEN 22 =>
						shift_out0 <= X352;
						shift_out1 <= X353;
						shift_out2 <= X354;
						shift_out3 <= X355;
						shift_out4 <= X356;
						shift_out5 <= X357;
						shift_out6 <= X358;
						shift_out7 <= X359;
						shift_out8 <= X360;
						shift_out9 <= X361;
						shift_out10 <= X362;
						shift_out11 <= X363;
						shift_out12 <= X364;
						shift_out13 <= X365;
						shift_out14 <= X366;
						shift_out15 <= X367;
						i <= i + 1;
					WHEN 23 =>
						shift_out0 <= X368;
						shift_out1 <= X369;
						shift_out2 <= X370;
						shift_out3 <= X371;
						shift_out4 <= X372;
						shift_out5 <= X373;
						shift_out6 <= X374;
						shift_out7 <= X375;
						shift_out8 <= X376;
						shift_out9 <= X377;
						shift_out10 <= X378;
						shift_out11 <= X379;
						shift_out12 <= X380;
						shift_out13 <= X381;
						shift_out14 <= X382;
						shift_out15 <= X383;
						i <= i + 1;
					WHEN 24 =>
						shift_out0 <= X384;
						shift_out1 <= X385;
						shift_out2 <= X386;
						shift_out3 <= X387;
						shift_out4 <= X388;
						shift_out5 <= X389;
						shift_out6 <= X390;
						shift_out7 <= X391;
						shift_out8 <= X392;
						shift_out9 <= X393;
						shift_out10 <= X394;
						shift_out11 <= X395;
						shift_out12 <= X396;
						shift_out13 <= X397;
						shift_out14 <= X398;
						shift_out15 <= X399;
						i <= i + 1;
					WHEN 25 =>
						shift_out0 <= X400;
						shift_out1 <= X401;
						shift_out2 <= X402;
						shift_out3 <= X403;
						shift_out4 <= X404;
						shift_out5 <= X405;
						shift_out6 <= X406;
						shift_out7 <= X407;
						shift_out8 <= X408;
						shift_out9 <= X409;
						shift_out10 <= X410;
						shift_out11 <= X411;
						shift_out12 <= X412;
						shift_out13 <= X413;
						shift_out14 <= X414;
						shift_out15 <= X415;
						i <= i + 1;
					WHEN 26 =>
						shift_out0 <= X416;
						shift_out1 <= X417;
						shift_out2 <= X418;
						shift_out3 <= X419;
						shift_out4 <= X420;
						shift_out5 <= X421;
						shift_out6 <= X422;
						shift_out7 <= X423;
						shift_out8 <= X424;
						shift_out9 <= X425;
						shift_out10 <= X426;
						shift_out11 <= X427;
						shift_out12 <= X428;
						shift_out13 <= X429;
						shift_out14 <= X430;
						shift_out15 <= X431;
						i <= i + 1;
					WHEN 27 =>
						shift_out0 <= X432;
						shift_out1 <= X433;
						shift_out2 <= X434;
						shift_out3 <= X435;
						shift_out4 <= X436;
						shift_out5 <= X437;
						shift_out6 <= X438;
						shift_out7 <= X439;
						shift_out8 <= X440;
						shift_out9 <= X441;
						shift_out10 <= X442;
						shift_out11 <= X443;
						shift_out12 <= X444;
						shift_out13 <= X445;
						shift_out14 <= X446;
						shift_out15 <= X447;
						i <= i + 1;
					WHEN 28 =>
						shift_out0 <= X448;
						shift_out1 <= X449;
						shift_out2 <= X450;
						shift_out3 <= X451;
						shift_out4 <= X452;
						shift_out5 <= X453;
						shift_out6 <= X454;
						shift_out7 <= X455;
						shift_out8 <= X456;
						shift_out9 <= X457;
						shift_out10 <= X458;
						shift_out11 <= X459;
						shift_out12 <= X460;
						shift_out13 <= X461;
						shift_out14 <= X462;
						shift_out15 <= X463;
						i <= i + 1;
					WHEN 29 =>
						shift_out0 <= X464;
						shift_out1 <= X465;
						shift_out2 <= X466;
						shift_out3 <= X467;
						shift_out4 <= X468;
						shift_out5 <= X469;
						shift_out6 <= X470;
						shift_out7 <= X471;
						shift_out8 <= X472;
						shift_out9 <= X473;
						shift_out10 <= X474;
						shift_out11 <= X475;
						shift_out12 <= X476;
						shift_out13 <= X477;
						shift_out14 <= X478;
						shift_out15 <= X479;
						i <= i + 1;
					WHEN 30 =>
						shift_out0 <= X480;
						shift_out1 <= X481;
						shift_out2 <= X482;
						shift_out3 <= X483;
						shift_out4 <= X484;
						shift_out5 <= X485;
						shift_out6 <= X486;
						shift_out7 <= X487;
						shift_out8 <= X488;
						shift_out9 <= X489;
						shift_out10 <= X490;
						shift_out11 <= X491;
						shift_out12 <= X492;
						shift_out13 <= X493;
						shift_out14 <= X494;
						shift_out15 <= X495;
						i <= i + 1;
					WHEN 31 =>
						shift_out0 <= X496;
						shift_out1 <= X497;
						shift_out2 <= X498;
						shift_out3 <= X499;
						shift_out4 <= X500;
						shift_out5 <= X501;
						shift_out6 <= X502;
						shift_out7 <= X503;
						shift_out8 <= X504;
						shift_out9 <= X505;
						shift_out10 <= X506;
						shift_out11 <= X507;
						shift_out12 <= X508;
						shift_out13 <= X509;
						shift_out14 <= X510;
						shift_out15 <= X511;
						i <= i + 1;
					WHEN 32 =>
						shift_out0 <= X512;
						shift_out1 <= X513;
						shift_out2 <= X514;
						shift_out3 <= X515;
						shift_out4 <= X516;
						shift_out5 <= X517;
						shift_out6 <= X518;
						shift_out7 <= X519;
						shift_out8 <= X520;
						shift_out9 <= X521;
						shift_out10 <= X522;
						shift_out11 <= X523;
						shift_out12 <= X524;
						shift_out13 <= X525;
						shift_out14 <= X526;
						shift_out15 <= X527;
						i <= i + 1;
					WHEN 33 =>
						shift_out0 <= X528;
						shift_out1 <= X529;
						shift_out2 <= X530;
						shift_out3 <= X531;
						shift_out4 <= X532;
						shift_out5 <= X533;
						shift_out6 <= X534;
						shift_out7 <= X535;
						shift_out8 <= X536;
						shift_out9 <= X537;
						shift_out10 <= X538;
						shift_out11 <= X539;
						shift_out12 <= X540;
						shift_out13 <= X541;
						shift_out14 <= X542;
						shift_out15 <= X543;
						i <= i + 1;
					WHEN 34 =>
						shift_out0 <= X544;
						shift_out1 <= X545;
						shift_out2 <= X546;
						shift_out3 <= X547;
						shift_out4 <= X548;
						shift_out5 <= X549;
						shift_out6 <= X550;
						shift_out7 <= X551;
						shift_out8 <= X552;
						shift_out9 <= X553;
						shift_out10 <= X554;
						shift_out11 <= X555;
						shift_out12 <= X556;
						shift_out13 <= X557;
						shift_out14 <= X558;
						shift_out15 <= X559;
						i <= i + 1;
					WHEN 35 =>
						shift_out0 <= X560;
						shift_out1 <= X561;
						shift_out2 <= X562;
						shift_out3 <= X563;
						shift_out4 <= X564;
						shift_out5 <= X565;
						shift_out6 <= X566;
						shift_out7 <= X567;
						shift_out8 <= X568;
						shift_out9 <= X569;
						shift_out10 <= X570;
						shift_out11 <= X571;
						shift_out12 <= X572;
						shift_out13 <= X573;
						shift_out14 <= X574;
						shift_out15 <= X575;
						i <= i + 1;
					WHEN 36 =>
						shift_out0 <= X576;
						shift_out1 <= X577;
						shift_out2 <= X578;
						shift_out3 <= X579;
						shift_out4 <= X580;
						shift_out5 <= X581;
						shift_out6 <= X582;
						shift_out7 <= X583;
						shift_out8 <= X584;
						shift_out9 <= X585;
						shift_out10 <= X586;
						shift_out11 <= X587;
						shift_out12 <= X588;
						shift_out13 <= X589;
						shift_out14 <= X590;
						shift_out15 <= X591;
						i <= i + 1;
					WHEN 37 =>
						shift_out0 <= X592;
						shift_out1 <= X593;
						shift_out2 <= X594;
						shift_out3 <= X595;
						shift_out4 <= X596;
						shift_out5 <= X597;
						shift_out6 <= X598;
						shift_out7 <= X599;
						shift_out8 <= X600;
						shift_out9 <= X601;
						shift_out10 <= X602;
						shift_out11 <= X603;
						shift_out12 <= X604;
						shift_out13 <= X605;
						shift_out14 <= X606;
						shift_out15 <= X607;
						i <= i + 1;
					WHEN 38 =>
						shift_out0 <= X608;
						shift_out1 <= X609;
						shift_out2 <= X610;
						shift_out3 <= X611;
						shift_out4 <= X612;
						shift_out5 <= X613;
						shift_out6 <= X614;
						shift_out7 <= X615;
						shift_out8 <= X616;
						shift_out9 <= X617;
						shift_out10 <= X618;
						shift_out11 <= X619;
						shift_out12 <= X620;
						shift_out13 <= X621;
						shift_out14 <= X622;
						shift_out15 <= X623;
						i <= i + 1;
					WHEN 39 =>
						shift_out0 <= X624;
						shift_out1 <= X625;
						shift_out2 <= X626;
						shift_out3 <= X627;
						shift_out4 <= X628;
						shift_out5 <= X629;
						shift_out6 <= X630;
						shift_out7 <= X631;
						shift_out8 <= X632;
						shift_out9 <= X633;
						shift_out10 <= X634;
						shift_out11 <= X635;
						shift_out12 <= X636;
						shift_out13 <= X637;
						shift_out14 <= X638;
						shift_out15 <= X639;
						i <= i + 1;
					WHEN 40 =>
						shift_out0 <= X640;
						shift_out1 <= X641;
						shift_out2 <= X642;
						shift_out3 <= X643;
						shift_out4 <= X644;
						shift_out5 <= X645;
						shift_out6 <= X646;
						shift_out7 <= X647;
						shift_out8 <= X648;
						shift_out9 <= X649;
						shift_out10 <= X650;
						shift_out11 <= X651;
						shift_out12 <= X652;
						shift_out13 <= X653;
						shift_out14 <= X654;
						shift_out15 <= X655;
						i <= i + 1;
					WHEN 41 =>
						shift_out0 <= X656;
						shift_out1 <= X657;
						shift_out2 <= X658;
						shift_out3 <= X659;
						shift_out4 <= X660;
						shift_out5 <= X661;
						shift_out6 <= X662;
						shift_out7 <= X663;
						shift_out8 <= X664;
						shift_out9 <= X665;
						shift_out10 <= X666;
						shift_out11 <= X667;
						shift_out12 <= X668;
						shift_out13 <= X669;
						shift_out14 <= X670;
						shift_out15 <= X671;
						i <= i + 1;
					WHEN 42 =>
						shift_out0 <= X672;
						shift_out1 <= X673;
						shift_out2 <= X674;
						shift_out3 <= X675;
						shift_out4 <= X676;
						shift_out5 <= X677;
						shift_out6 <= X678;
						shift_out7 <= X679;
						shift_out8 <= X680;
						shift_out9 <= X681;
						shift_out10 <= X682;
						shift_out11 <= X683;
						shift_out12 <= X684;
						shift_out13 <= X685;
						shift_out14 <= X686;
						shift_out15 <= X687;
						i <= i + 1;
					WHEN 43 =>
						shift_out0 <= X688;
						shift_out1 <= X689;
						shift_out2 <= X690;
						shift_out3 <= X691;
						shift_out4 <= X692;
						shift_out5 <= X693;
						shift_out6 <= X694;
						shift_out7 <= X695;
						shift_out8 <= X696;
						shift_out9 <= X697;
						shift_out10 <= X698;
						shift_out11 <= X699;
						shift_out12 <= X700;
						shift_out13 <= X701;
						shift_out14 <= X702;
						shift_out15 <= X703;
						i <= i + 1;
					WHEN 44 =>
						shift_out0 <= X704;
						shift_out1 <= X705;
						shift_out2 <= X706;
						shift_out3 <= X707;
						shift_out4 <= X708;
						shift_out5 <= X709;
						shift_out6 <= X710;
						shift_out7 <= X711;
						shift_out8 <= X712;
						shift_out9 <= X713;
						shift_out10 <= X714;
						shift_out11 <= X715;
						shift_out12 <= X716;
						shift_out13 <= X717;
						shift_out14 <= X718;
						shift_out15 <= X719;
						i <= i + 1;
					WHEN 45 =>
						shift_out0 <= X720;
						shift_out1 <= X721;
						shift_out2 <= X722;
						shift_out3 <= X723;
						shift_out4 <= X724;
						shift_out5 <= X725;
						shift_out6 <= X726;
						shift_out7 <= X727;
						shift_out8 <= X728;
						shift_out9 <= X729;
						shift_out10 <= X730;
						shift_out11 <= X731;
						shift_out12 <= X732;
						shift_out13 <= X733;
						shift_out14 <= X734;
						shift_out15 <= X735;
						i <= i + 1;
					WHEN 46 =>
						shift_out0 <= X736;
						shift_out1 <= X737;
						shift_out2 <= X738;
						shift_out3 <= X739;
						shift_out4 <= X740;
						shift_out5 <= X741;
						shift_out6 <= X742;
						shift_out7 <= X743;
						shift_out8 <= X744;
						shift_out9 <= X745;
						shift_out10 <= X746;
						shift_out11 <= X747;
						shift_out12 <= X748;
						shift_out13 <= X749;
						shift_out14 <= X750;
						shift_out15 <= X751;
						i <= i + 1;
					WHEN 47 =>
						shift_out0 <= X752;
						shift_out1 <= X753;
						shift_out2 <= X754;
						shift_out3 <= X755;
						shift_out4 <= X756;
						shift_out5 <= X757;
						shift_out6 <= X758;
						shift_out7 <= X759;
						shift_out8 <= X760;
						shift_out9 <= X761;
						shift_out10 <= X762;
						shift_out11 <= X763;
						shift_out12 <= X764;
						shift_out13 <= X765;
						shift_out14 <= X766;
						shift_out15 <= X767;
						i <= i + 1;
					WHEN 48 =>
						shift_out0 <= X768;
						shift_out1 <= X769;
						shift_out2 <= X770;
						shift_out3 <= X771;
						shift_out4 <= X772;
						shift_out5 <= X773;
						shift_out6 <= X774;
						shift_out7 <= X775;
						shift_out8 <= X776;
						shift_out9 <= X777;
						shift_out10 <= X778;
						shift_out11 <= X779;
						shift_out12 <= X780;
						shift_out13 <= X781;
						shift_out14 <= X782;
						shift_out15 <= X783;
						i <= i + 1;
					WHEN 49 =>
						shift_out0 <= X784;
						shift_out1 <= X785;
						shift_out2 <= X786;
						shift_out3 <= X787;
						shift_out4 <= X788;
						shift_out5 <= X789;
						shift_out6 <= X790;
						shift_out7 <= X791;
						shift_out8 <= X792;
						shift_out9 <= X793;
						shift_out10 <= X794;
						shift_out11 <= X795;
						shift_out12 <= X796;
						shift_out13 <= X797;
						shift_out14 <= X798;
						shift_out15 <= X799;
						i <= i + 1;
					WHEN 50 =>
						shift_out0 <= X800;
						shift_out1 <= X801;
						shift_out2 <= X802;
						shift_out3 <= X803;
						shift_out4 <= X804;
						shift_out5 <= X805;
						shift_out6 <= X806;
						shift_out7 <= X807;
						shift_out8 <= X808;
						shift_out9 <= X809;
						shift_out10 <= X810;
						shift_out11 <= X811;
						shift_out12 <= X812;
						shift_out13 <= X813;
						shift_out14 <= X814;
						shift_out15 <= X815;
						i <= i + 1;
					WHEN 51 =>
						shift_out0 <= X816;
						shift_out1 <= X817;
						shift_out2 <= X818;
						shift_out3 <= X819;
						shift_out4 <= X820;
						shift_out5 <= X821;
						shift_out6 <= X822;
						shift_out7 <= X823;
						shift_out8 <= X824;
						shift_out9 <= X825;
						shift_out10 <= X826;
						shift_out11 <= X827;
						shift_out12 <= X828;
						shift_out13 <= X829;
						shift_out14 <= X830;
						shift_out15 <= X831;
						i <= i + 1;
					WHEN 52 =>
						shift_out0 <= X832;
						shift_out1 <= X833;
						shift_out2 <= X834;
						shift_out3 <= X835;
						shift_out4 <= X836;
						shift_out5 <= X837;
						shift_out6 <= X838;
						shift_out7 <= X839;
						shift_out8 <= X840;
						shift_out9 <= X841;
						shift_out10 <= X842;
						shift_out11 <= X843;
						shift_out12 <= X844;
						shift_out13 <= X845;
						shift_out14 <= X846;
						shift_out15 <= X847;
						i <= i + 1;
					WHEN 53 =>
						shift_out0 <= X848;
						shift_out1 <= X849;
						shift_out2 <= X850;
						shift_out3 <= X851;
						shift_out4 <= X852;
						shift_out5 <= X853;
						shift_out6 <= X854;
						shift_out7 <= X855;
						shift_out8 <= X856;
						shift_out9 <= X857;
						shift_out10 <= X858;
						shift_out11 <= X859;
						shift_out12 <= X860;
						shift_out13 <= X861;
						shift_out14 <= X862;
						shift_out15 <= X863;
						i <= i + 1;
					WHEN 54 =>
						shift_out0 <= X864;
						shift_out1 <= X865;
						shift_out2 <= X866;
						shift_out3 <= X867;
						shift_out4 <= X868;
						shift_out5 <= X869;
						shift_out6 <= X870;
						shift_out7 <= X871;
						shift_out8 <= X872;
						shift_out9 <= X873;
						shift_out10 <= X874;
						shift_out11 <= X875;
						shift_out12 <= X876;
						shift_out13 <= X877;
						shift_out14 <= X878;
						shift_out15 <= X879;
						i <= i + 1;
					WHEN 55 =>
						shift_out0 <= X880;
						shift_out1 <= X881;
						shift_out2 <= X882;
						shift_out3 <= X883;
						shift_out4 <= X884;
						shift_out5 <= X885;
						shift_out6 <= X886;
						shift_out7 <= X887;
						shift_out8 <= X888;
						shift_out9 <= X889;
						shift_out10 <= X890;
						shift_out11 <= X891;
						shift_out12 <= X892;
						shift_out13 <= X893;
						shift_out14 <= X894;
						shift_out15 <= X895;
						i <= i + 1;
					WHEN 56 =>
						shift_out0 <= X896;
						shift_out1 <= X897;
						shift_out2 <= X898;
						shift_out3 <= X899;
						shift_out4 <= X900;
						shift_out5 <= X901;
						shift_out6 <= X902;
						shift_out7 <= X903;
						shift_out8 <= X904;
						shift_out9 <= X905;
						shift_out10 <= X906;
						shift_out11 <= X907;
						shift_out12 <= X908;
						shift_out13 <= X909;
						shift_out14 <= X910;
						shift_out15 <= X911;
						i <= i + 1;
					WHEN 57 =>
						shift_out0 <= X912;
						shift_out1 <= X913;
						shift_out2 <= X914;
						shift_out3 <= X915;
						shift_out4 <= X916;
						shift_out5 <= X917;
						shift_out6 <= X918;
						shift_out7 <= X919;
						shift_out8 <= X920;
						shift_out9 <= X921;
						shift_out10 <= X922;
						shift_out11 <= X923;
						shift_out12 <= X924;
						shift_out13 <= X925;
						shift_out14 <= X926;
						shift_out15 <= X927;
						i <= i + 1;
					WHEN 58 =>
						shift_out0 <= X928;
						shift_out1 <= X929;
						shift_out2 <= X930;
						shift_out3 <= X931;
						shift_out4 <= X932;
						shift_out5 <= X933;
						shift_out6 <= X934;
						shift_out7 <= X935;
						shift_out8 <= X936;
						shift_out9 <= X937;
						shift_out10 <= X938;
						shift_out11 <= X939;
						shift_out12 <= X940;
						shift_out13 <= X941;
						shift_out14 <= X942;
						shift_out15 <= X943;
						i <= i + 1;
					WHEN 59 =>
						shift_out0 <= X944;
						shift_out1 <= X945;
						shift_out2 <= X946;
						shift_out3 <= X947;
						shift_out4 <= X948;
						shift_out5 <= X949;
						shift_out6 <= X950;
						shift_out7 <= X951;
						shift_out8 <= X952;
						shift_out9 <= X953;
						shift_out10 <= X954;
						shift_out11 <= X955;
						shift_out12 <= X956;
						shift_out13 <= X957;
						shift_out14 <= X958;
						shift_out15 <= X959;
						i <= i + 1;
					WHEN 60 =>
						shift_out0 <= X960;
						shift_out1 <= X961;
						shift_out2 <= X962;
						shift_out3 <= X963;
						shift_out4 <= X964;
						shift_out5 <= X965;
						shift_out6 <= X966;
						shift_out7 <= X967;
						shift_out8 <= X968;
						shift_out9 <= X969;
						shift_out10 <= X970;
						shift_out11 <= X971;
						shift_out12 <= X972;
						shift_out13 <= X973;
						shift_out14 <= X974;
						shift_out15 <= X975;
						i <= i + 1;
					WHEN 61 =>
						shift_out0 <= X976;
						shift_out1 <= X977;
						shift_out2 <= X978;
						shift_out3 <= X979;
						shift_out4 <= X980;
						shift_out5 <= X981;
						shift_out6 <= X982;
						shift_out7 <= X983;
						shift_out8 <= X984;
						shift_out9 <= X985;
						shift_out10 <= X986;
						shift_out11 <= X987;
						shift_out12 <= X988;
						shift_out13 <= X989;
						shift_out14 <= X990;
						shift_out15 <= X991;
						i <= i + 1;
					WHEN 62 =>
						shift_out0 <= X992;
						shift_out1 <= X993;
						shift_out2 <= X994;
						shift_out3 <= X995;
						shift_out4 <= X996;
						shift_out5 <= X997;
						shift_out6 <= X998;
						shift_out7 <= X999;
						shift_out8 <= X1000;
						shift_out9 <= X1001;
						shift_out10 <= X1002;
						shift_out11 <= X1003;
						shift_out12 <= X1004;
						shift_out13 <= X1005;
						shift_out14 <= X1006;
						shift_out15 <= X1007;
						i <= i + 1;
					WHEN 63 =>
						shift_out0 <= X1008;
						shift_out1 <= X1009;
						shift_out2 <= X1010;
						shift_out3 <= X1011;
						shift_out4 <= X1012;
						shift_out5 <= X1013;
						shift_out6 <= X1014;
						shift_out7 <= X1015;
						shift_out8 <= X1016;
						shift_out9 <= X1017;
						shift_out10 <= X1018;
						shift_out11 <= X1019;
						shift_out12 <= X1020;
						shift_out13 <= X1021;
						shift_out14 <= X1022;
						shift_out15 <= X1023;
						i <= i + 1;
					WHEN 64 =>
						shift_out0 <= X1024;
						shift_out1 <= X1025;
						shift_out2 <= X1026;
						shift_out3 <= X1027;
						shift_out4 <= X1028;
						shift_out5 <= X1029;
						shift_out6 <= X1030;
						shift_out7 <= X1031;
						shift_out8 <= X1032;
						shift_out9 <= X1033;
						shift_out10 <= X1034;
						shift_out11 <= X1035;
						shift_out12 <= X1036;
						shift_out13 <= X1037;
						shift_out14 <= X1038;
						shift_out15 <= X1039;
						i <= i + 1;
					WHEN 65 =>
						shift_out0 <= X1040;
						shift_out1 <= X1041;
						shift_out2 <= X1042;
						shift_out3 <= X1043;
						shift_out4 <= X1044;
						shift_out5 <= X1045;
						shift_out6 <= X1046;
						shift_out7 <= X1047;
						shift_out8 <= X1048;
						shift_out9 <= X1049;
						shift_out10 <= X1050;
						shift_out11 <= X1051;
						shift_out12 <= X1052;
						shift_out13 <= X1053;
						shift_out14 <= X1054;
						shift_out15 <= X1055;
						i <= i + 1;
					WHEN 66 =>
						shift_out0 <= X1056;
						shift_out1 <= X1057;
						shift_out2 <= X1058;
						shift_out3 <= X1059;
						shift_out4 <= X1060;
						shift_out5 <= X1061;
						shift_out6 <= X1062;
						shift_out7 <= X1063;
						shift_out8 <= X1064;
						shift_out9 <= X1065;
						shift_out10 <= X1066;
						shift_out11 <= X1067;
						shift_out12 <= X1068;
						shift_out13 <= X1069;
						shift_out14 <= X1070;
						shift_out15 <= X1071;
						i <= i + 1;
					WHEN 67 =>
						shift_out0 <= X1072;
						shift_out1 <= X1073;
						shift_out2 <= X1074;
						shift_out3 <= X1075;
						shift_out4 <= X1076;
						shift_out5 <= X1077;
						shift_out6 <= X1078;
						shift_out7 <= X1079;
						shift_out8 <= X1080;
						shift_out9 <= X1081;
						shift_out10 <= X1082;
						shift_out11 <= X1083;
						shift_out12 <= X1084;
						shift_out13 <= X1085;
						shift_out14 <= X1086;
						shift_out15 <= X1087;
						i <= i + 1;
					WHEN 68 =>
						shift_out0 <= X1088;
						shift_out1 <= X1089;
						shift_out2 <= X1090;
						shift_out3 <= X1091;
						shift_out4 <= X1092;
						shift_out5 <= X1093;
						shift_out6 <= X1094;
						shift_out7 <= X1095;
						shift_out8 <= X1096;
						shift_out9 <= X1097;
						shift_out10 <= X1098;
						shift_out11 <= X1099;
						shift_out12 <= X1100;
						shift_out13 <= X1101;
						shift_out14 <= X1102;
						shift_out15 <= X1103;
						i <= i + 1;
					WHEN 69 =>
						shift_out0 <= X1104;
						shift_out1 <= X1105;
						shift_out2 <= X1106;
						shift_out3 <= X1107;
						shift_out4 <= X1108;
						shift_out5 <= X1109;
						shift_out6 <= X1110;
						shift_out7 <= X1111;
						shift_out8 <= X1112;
						shift_out9 <= X1113;
						shift_out10 <= X1114;
						shift_out11 <= X1115;
						shift_out12 <= X1116;
						shift_out13 <= X1117;
						shift_out14 <= X1118;
						shift_out15 <= X1119;
						i <= i + 1;
					WHEN 70 =>
						shift_out0 <= X1120;
						shift_out1 <= X1121;
						shift_out2 <= X1122;
						shift_out3 <= X1123;
						shift_out4 <= X1124;
						shift_out5 <= X1125;
						shift_out6 <= X1126;
						shift_out7 <= X1127;
						shift_out8 <= X1128;
						shift_out9 <= X1129;
						shift_out10 <= X1130;
						shift_out11 <= X1131;
						shift_out12 <= X1132;
						shift_out13 <= X1133;
						shift_out14 <= X1134;
						shift_out15 <= X1135;
						i <= i + 1;
					WHEN 71 =>
						shift_out0 <= X1136;
						shift_out1 <= X1137;
						shift_out2 <= X1138;
						shift_out3 <= X1139;
						shift_out4 <= X1140;
						shift_out5 <= X1141;
						shift_out6 <= X1142;
						shift_out7 <= X1143;
						shift_out8 <= X1144;
						shift_out9 <= X1145;
						shift_out10 <= X1146;
						shift_out11 <= X1147;
						shift_out12 <= X1148;
						shift_out13 <= X1149;
						shift_out14 <= X1150;
						shift_out15 <= X1151;
						i <= i + 1;
					WHEN 72 =>
						shift_out0 <= X1152;
						shift_out1 <= X1153;
						shift_out2 <= X1154;
						shift_out3 <= X1155;
						shift_out4 <= X1156;
						shift_out5 <= X1157;
						shift_out6 <= X1158;
						shift_out7 <= X1159;
						shift_out8 <= X1160;
						shift_out9 <= X1161;
						shift_out10 <= X1162;
						shift_out11 <= X1163;
						shift_out12 <= X1164;
						shift_out13 <= X1165;
						shift_out14 <= X1166;
						shift_out15 <= X1167;
						i <= i + 1;
					WHEN 73 =>
						shift_out0 <= X1168;
						shift_out1 <= X1169;
						shift_out2 <= X1170;
						shift_out3 <= X1171;
						shift_out4 <= X1172;
						shift_out5 <= X1173;
						shift_out6 <= X1174;
						shift_out7 <= X1175;
						shift_out8 <= X1176;
						shift_out9 <= X1177;
						shift_out10 <= X1178;
						shift_out11 <= X1179;
						shift_out12 <= X1180;
						shift_out13 <= X1181;
						shift_out14 <= X1182;
						shift_out15 <= X1183;
						i <= i + 1;
					WHEN 74 =>
						shift_out0 <= X1184;
						shift_out1 <= X1185;
						shift_out2 <= X1186;
						shift_out3 <= X1187;
						shift_out4 <= X1188;
						shift_out5 <= X1189;
						shift_out6 <= X1190;
						shift_out7 <= X1191;
						shift_out8 <= X1192;
						shift_out9 <= X1193;
						shift_out10 <= X1194;
						shift_out11 <= X1195;
						shift_out12 <= X1196;
						shift_out13 <= X1197;
						shift_out14 <= X1198;
						shift_out15 <= X1199;
						i <= i + 1;
					WHEN 75 =>
						shift_out0 <= X1200;
						shift_out1 <= X1201;
						shift_out2 <= X1202;
						shift_out3 <= X1203;
						shift_out4 <= X1204;
						shift_out5 <= X1205;
						shift_out6 <= X1206;
						shift_out7 <= X1207;
						shift_out8 <= X1208;
						shift_out9 <= X1209;
						shift_out10 <= X1210;
						shift_out11 <= X1211;
						shift_out12 <= X1212;
						shift_out13 <= X1213;
						shift_out14 <= X1214;
						shift_out15 <= X1215;
						i <= i + 1;
					WHEN 76 =>
						shift_out0 <= X1216;
						shift_out1 <= X1217;
						shift_out2 <= X1218;
						shift_out3 <= X1219;
						shift_out4 <= X1220;
						shift_out5 <= X1221;
						shift_out6 <= X1222;
						shift_out7 <= X1223;
						shift_out8 <= X1224;
						shift_out9 <= X1225;
						shift_out10 <= X1226;
						shift_out11 <= X1227;
						shift_out12 <= X1228;
						shift_out13 <= X1229;
						shift_out14 <= X1230;
						shift_out15 <= X1231;
						i <= i + 1;
					WHEN 77 =>
						shift_out0 <= X1232;
						shift_out1 <= X1233;
						shift_out2 <= X1234;
						shift_out3 <= X1235;
						shift_out4 <= X1236;
						shift_out5 <= X1237;
						shift_out6 <= X1238;
						shift_out7 <= X1239;
						shift_out8 <= X1240;
						shift_out9 <= X1241;
						shift_out10 <= X1242;
						shift_out11 <= X1243;
						shift_out12 <= X1244;
						shift_out13 <= X1245;
						shift_out14 <= X1246;
						shift_out15 <= X1247;
						i <= i + 1;
					WHEN 78 =>
						shift_out0 <= X1248;
						shift_out1 <= X1249;
						shift_out2 <= X1250;
						shift_out3 <= X1251;
						shift_out4 <= X1252;
						shift_out5 <= X1253;
						shift_out6 <= X1254;
						shift_out7 <= X1255;
						shift_out8 <= X1256;
						shift_out9 <= X1257;
						shift_out10 <= X1258;
						shift_out11 <= X1259;
						shift_out12 <= X1260;
						shift_out13 <= X1261;
						shift_out14 <= X1262;
						shift_out15 <= X1263;
						i <= i + 1;
					WHEN 79 =>
						shift_out0 <= X1264;
						shift_out1 <= X1265;
						shift_out2 <= X1266;
						shift_out3 <= X1267;
						shift_out4 <= X1268;
						shift_out5 <= X1269;
						shift_out6 <= X1270;
						shift_out7 <= X1271;
						shift_out8 <= X1272;
						shift_out9 <= X1273;
						shift_out10 <= X1274;
						shift_out11 <= X1275;
						shift_out12 <= X1276;
						shift_out13 <= X1277;
						shift_out14 <= X1278;
						shift_out15 <= X1279;
						i <= i + 1;
					WHEN 80 =>
						shift_out0 <= X1280;
						shift_out1 <= X1281;
						shift_out2 <= X1282;
						shift_out3 <= X1283;
						shift_out4 <= X1284;
						shift_out5 <= X1285;
						shift_out6 <= X1286;
						shift_out7 <= X1287;
						shift_out8 <= X1288;
						shift_out9 <= X1289;
						shift_out10 <= X1290;
						shift_out11 <= X1291;
						shift_out12 <= X1292;
						shift_out13 <= X1293;
						shift_out14 <= X1294;
						shift_out15 <= X1295;
						i <= i + 1;
					WHEN 81 =>
						shift_out0 <= X1296;
						shift_out1 <= X1297;
						shift_out2 <= X1298;
						shift_out3 <= X1299;
						shift_out4 <= X1300;
						shift_out5 <= X1301;
						shift_out6 <= X1302;
						shift_out7 <= X1303;
						shift_out8 <= X1304;
						shift_out9 <= X1305;
						shift_out10 <= X1306;
						shift_out11 <= X1307;
						shift_out12 <= X1308;
						shift_out13 <= X1309;
						shift_out14 <= X1310;
						shift_out15 <= X1311;
						i <= i + 1;
					WHEN 82 =>
						shift_out0 <= X1312;
						shift_out1 <= X1313;
						shift_out2 <= X1314;
						shift_out3 <= X1315;
						shift_out4 <= X1316;
						shift_out5 <= X1317;
						shift_out6 <= X1318;
						shift_out7 <= X1319;
						shift_out8 <= X1320;
						shift_out9 <= X1321;
						shift_out10 <= X1322;
						shift_out11 <= X1323;
						shift_out12 <= X1324;
						shift_out13 <= X1325;
						shift_out14 <= X1326;
						shift_out15 <= X1327;
						i <= i + 1;
					WHEN 83 =>
						shift_out0 <= X1328;
						shift_out1 <= X1329;
						shift_out2 <= X1330;
						shift_out3 <= X1331;
						shift_out4 <= X1332;
						shift_out5 <= X1333;
						shift_out6 <= X1334;
						shift_out7 <= X1335;
						shift_out8 <= X1336;
						shift_out9 <= X1337;
						shift_out10 <= X1338;
						shift_out11 <= X1339;
						shift_out12 <= X1340;
						shift_out13 <= X1341;
						shift_out14 <= X1342;
						shift_out15 <= X1343;
						i <= i + 1;
					WHEN 84 =>
						shift_out0 <= X1344;
						shift_out1 <= X1345;
						shift_out2 <= X1346;
						shift_out3 <= X1347;
						shift_out4 <= X1348;
						shift_out5 <= X1349;
						shift_out6 <= X1350;
						shift_out7 <= X1351;
						shift_out8 <= X1352;
						shift_out9 <= X1353;
						shift_out10 <= X1354;
						shift_out11 <= X1355;
						shift_out12 <= X1356;
						shift_out13 <= X1357;
						shift_out14 <= X1358;
						shift_out15 <= X1359;
						i <= i + 1;
					WHEN 85 =>
						shift_out0 <= X1360;
						shift_out1 <= X1361;
						shift_out2 <= X1362;
						shift_out3 <= X1363;
						shift_out4 <= X1364;
						shift_out5 <= X1365;
						shift_out6 <= X1366;
						shift_out7 <= X1367;
						shift_out8 <= X1368;
						shift_out9 <= X1369;
						shift_out10 <= X1370;
						shift_out11 <= X1371;
						shift_out12 <= X1372;
						shift_out13 <= X1373;
						shift_out14 <= X1374;
						shift_out15 <= X1375;
						i <= i + 1;
					WHEN 86 =>
						shift_out0 <= X1376;
						shift_out1 <= X1377;
						shift_out2 <= X1378;
						shift_out3 <= X1379;
						shift_out4 <= X1380;
						shift_out5 <= X1381;
						shift_out6 <= X1382;
						shift_out7 <= X1383;
						shift_out8 <= X1384;
						shift_out9 <= X1385;
						shift_out10 <= X1386;
						shift_out11 <= X1387;
						shift_out12 <= X1388;
						shift_out13 <= X1389;
						shift_out14 <= X1390;
						shift_out15 <= X1391;
						i <= i + 1;
					WHEN 87 =>
						shift_out0 <= X1392;
						shift_out1 <= X1393;
						shift_out2 <= X1394;
						shift_out3 <= X1395;
						shift_out4 <= X1396;
						shift_out5 <= X1397;
						shift_out6 <= X1398;
						shift_out7 <= X1399;
						shift_out8 <= X1400;
						shift_out9 <= X1401;
						shift_out10 <= X1402;
						shift_out11 <= X1403;
						shift_out12 <= X1404;
						shift_out13 <= X1405;
						shift_out14 <= X1406;
						shift_out15 <= X1407;
						i <= i + 1;
					WHEN 88 =>
						shift_out0 <= X1408;
						shift_out1 <= X1409;
						shift_out2 <= X1410;
						shift_out3 <= X1411;
						shift_out4 <= X1412;
						shift_out5 <= X1413;
						shift_out6 <= X1414;
						shift_out7 <= X1415;
						shift_out8 <= X1416;
						shift_out9 <= X1417;
						shift_out10 <= X1418;
						shift_out11 <= X1419;
						shift_out12 <= X1420;
						shift_out13 <= X1421;
						shift_out14 <= X1422;
						shift_out15 <= X1423;
						i <= i + 1;
					WHEN 89 =>
						shift_out0 <= X1424;
						shift_out1 <= X1425;
						shift_out2 <= X1426;
						shift_out3 <= X1427;
						shift_out4 <= X1428;
						shift_out5 <= X1429;
						shift_out6 <= X1430;
						shift_out7 <= X1431;
						shift_out8 <= X1432;
						shift_out9 <= X1433;
						shift_out10 <= X1434;
						shift_out11 <= X1435;
						shift_out12 <= X1436;
						shift_out13 <= X1437;
						shift_out14 <= X1438;
						shift_out15 <= X1439;
						i <= i + 1;
					WHEN 90 =>
						shift_out0 <= X1440;
						shift_out1 <= X1441;
						shift_out2 <= X1442;
						shift_out3 <= X1443;
						shift_out4 <= X1444;
						shift_out5 <= X1445;
						shift_out6 <= X1446;
						shift_out7 <= X1447;
						shift_out8 <= X1448;
						shift_out9 <= X1449;
						shift_out10 <= X1450;
						shift_out11 <= X1451;
						shift_out12 <= X1452;
						shift_out13 <= X1453;
						shift_out14 <= X1454;
						shift_out15 <= X1455;
						i <= i + 1;
					WHEN 91 =>
						shift_out0 <= X1456;
						shift_out1 <= X1457;
						shift_out2 <= X1458;
						shift_out3 <= X1459;
						shift_out4 <= X1460;
						shift_out5 <= X1461;
						shift_out6 <= X1462;
						shift_out7 <= X1463;
						shift_out8 <= X1464;
						shift_out9 <= X1465;
						shift_out10 <= X1466;
						shift_out11 <= X1467;
						shift_out12 <= X1468;
						shift_out13 <= X1469;
						shift_out14 <= X1470;
						shift_out15 <= X1471;
						i <= i + 1;
					WHEN 92 =>
						shift_out0 <= X1472;
						shift_out1 <= X1473;
						shift_out2 <= X1474;
						shift_out3 <= X1475;
						shift_out4 <= X1476;
						shift_out5 <= X1477;
						shift_out6 <= X1478;
						shift_out7 <= X1479;
						shift_out8 <= X1480;
						shift_out9 <= X1481;
						shift_out10 <= X1482;
						shift_out11 <= X1483;
						shift_out12 <= X1484;
						shift_out13 <= X1485;
						shift_out14 <= X1486;
						shift_out15 <= X1487;
						i <= i + 1;
					WHEN 93 =>
						shift_out0 <= X1488;
						shift_out1 <= X1489;
						shift_out2 <= X1490;
						shift_out3 <= X1491;
						shift_out4 <= X1492;
						shift_out5 <= X1493;
						shift_out6 <= X1494;
						shift_out7 <= X1495;
						shift_out8 <= X1496;
						shift_out9 <= X1497;
						shift_out10 <= X1498;
						shift_out11 <= X1499;
						shift_out12 <= X1500;
						shift_out13 <= X1501;
						shift_out14 <= X1502;
						shift_out15 <= X1503;
						i <= i + 1;
					WHEN 94 =>
						shift_out0 <= X1504;
						shift_out1 <= X1505;
						shift_out2 <= X1506;
						shift_out3 <= X1507;
						shift_out4 <= X1508;
						shift_out5 <= X1509;
						shift_out6 <= X1510;
						shift_out7 <= X1511;
						shift_out8 <= X1512;
						shift_out9 <= X1513;
						shift_out10 <= X1514;
						shift_out11 <= X1515;
						shift_out12 <= X1516;
						shift_out13 <= X1517;
						shift_out14 <= X1518;
						shift_out15 <= X1519;
						i <= i + 1;
					WHEN 95 =>
						shift_out0 <= X1520;
						shift_out1 <= X1521;
						shift_out2 <= X1522;
						shift_out3 <= X1523;
						shift_out4 <= X1524;
						shift_out5 <= X1525;
						shift_out6 <= X1526;
						shift_out7 <= X1527;
						shift_out8 <= X1528;
						shift_out9 <= X1529;
						shift_out10 <= X1530;
						shift_out11 <= X1531;
						shift_out12 <= X1532;
						shift_out13 <= X1533;
						shift_out14 <= X1534;
						shift_out15 <= X1535;
						i <= i + 1;
					WHEN 96 =>
						shift_out0 <= X1536;
						shift_out1 <= X1537;
						shift_out2 <= X1538;
						shift_out3 <= X1539;
						shift_out4 <= X1540;
						shift_out5 <= X1541;
						shift_out6 <= X1542;
						shift_out7 <= X1543;
						shift_out8 <= X1544;
						shift_out9 <= X1545;
						shift_out10 <= X1546;
						shift_out11 <= X1547;
						shift_out12 <= X1548;
						shift_out13 <= X1549;
						shift_out14 <= X1550;
						shift_out15 <= X1551;
						i <= i + 1;
					WHEN 97 =>
						shift_out0 <= X1552;
						shift_out1 <= X1553;
						shift_out2 <= X1554;
						shift_out3 <= X1555;
						shift_out4 <= X1556;
						shift_out5 <= X1557;
						shift_out6 <= X1558;
						shift_out7 <= X1559;
						shift_out8 <= X1560;
						shift_out9 <= X1561;
						shift_out10 <= X1562;
						shift_out11 <= X1563;
						shift_out12 <= X1564;
						shift_out13 <= X1565;
						shift_out14 <= X1566;
						shift_out15 <= X1567;
						i <= i + 1;
					WHEN 98 =>
						shift_out0 <= X1568;
						shift_out1 <= X1569;
						shift_out2 <= X1570;
						shift_out3 <= X1571;
						shift_out4 <= X1572;
						shift_out5 <= X1573;
						shift_out6 <= X1574;
						shift_out7 <= X1575;
						shift_out8 <= X1576;
						shift_out9 <= X1577;
						shift_out10 <= X1578;
						shift_out11 <= X1579;
						shift_out12 <= X1580;
						shift_out13 <= X1581;
						shift_out14 <= X1582;
						shift_out15 <= X1583;
						i <= i + 1;
					WHEN 99 =>
						shift_out0 <= X1584;
						shift_out1 <= X1585;
						shift_out2 <= X1586;
						shift_out3 <= X1587;
						shift_out4 <= X1588;
						shift_out5 <= X1589;
						shift_out6 <= X1590;
						shift_out7 <= X1591;
						shift_out8 <= X1592;
						shift_out9 <= X1593;
						shift_out10 <= X1594;
						shift_out11 <= X1595;
						shift_out12 <= X1596;
						shift_out13 <= X1597;
						shift_out14 <= X1598;
						shift_out15 <= X1599;
						i <= i + 1;
					WHEN 100 =>
						shift_out0 <= X1600;
						shift_out1 <= X1601;
						shift_out2 <= X1602;
						shift_out3 <= X1603;
						shift_out4 <= X1604;
						shift_out5 <= X1605;
						shift_out6 <= X1606;
						shift_out7 <= X1607;
						shift_out8 <= X1608;
						shift_out9 <= X1609;
						shift_out10 <= X1610;
						shift_out11 <= X1611;
						shift_out12 <= X1612;
						shift_out13 <= X1613;
						shift_out14 <= X1614;
						shift_out15 <= X1615;
						i <= i + 1;
					WHEN 101 =>
						shift_out0 <= X1616;
						shift_out1 <= X1617;
						shift_out2 <= X1618;
						shift_out3 <= X1619;
						shift_out4 <= X1620;
						shift_out5 <= X1621;
						shift_out6 <= X1622;
						shift_out7 <= X1623;
						shift_out8 <= X1624;
						shift_out9 <= X1625;
						shift_out10 <= X1626;
						shift_out11 <= X1627;
						shift_out12 <= X1628;
						shift_out13 <= X1629;
						shift_out14 <= X1630;
						shift_out15 <= X1631;
						i <= i + 1;
					WHEN 102 =>
						shift_out0 <= X1632;
						shift_out1 <= X1633;
						shift_out2 <= X1634;
						shift_out3 <= X1635;
						shift_out4 <= X1636;
						shift_out5 <= X1637;
						shift_out6 <= X1638;
						shift_out7 <= X1639;
						shift_out8 <= X1640;
						shift_out9 <= X1641;
						shift_out10 <= X1642;
						shift_out11 <= X1643;
						shift_out12 <= X1644;
						shift_out13 <= X1645;
						shift_out14 <= X1646;
						shift_out15 <= X1647;
						i <= i + 1;
					WHEN 103 =>
						shift_out0 <= X1648;
						shift_out1 <= X1649;
						shift_out2 <= X1650;
						shift_out3 <= X1651;
						shift_out4 <= X1652;
						shift_out5 <= X1653;
						shift_out6 <= X1654;
						shift_out7 <= X1655;
						shift_out8 <= X1656;
						shift_out9 <= X1657;
						shift_out10 <= X1658;
						shift_out11 <= X1659;
						shift_out12 <= X1660;
						shift_out13 <= X1661;
						shift_out14 <= X1662;
						shift_out15 <= X1663;
						i <= i + 1;
					WHEN 104 =>
						shift_out0 <= X1664;
						shift_out1 <= X1665;
						shift_out2 <= X1666;
						shift_out3 <= X1667;
						shift_out4 <= X1668;
						shift_out5 <= X1669;
						shift_out6 <= X1670;
						shift_out7 <= X1671;
						shift_out8 <= X1672;
						shift_out9 <= X1673;
						shift_out10 <= X1674;
						shift_out11 <= X1675;
						shift_out12 <= X1676;
						shift_out13 <= X1677;
						shift_out14 <= X1678;
						shift_out15 <= X1679;
						i <= i + 1;
					WHEN 105 =>
						shift_out0 <= X1680;
						shift_out1 <= X1681;
						shift_out2 <= X1682;
						shift_out3 <= X1683;
						shift_out4 <= X1684;
						shift_out5 <= X1685;
						shift_out6 <= X1686;
						shift_out7 <= X1687;
						shift_out8 <= X1688;
						shift_out9 <= X1689;
						shift_out10 <= X1690;
						shift_out11 <= X1691;
						shift_out12 <= X1692;
						shift_out13 <= X1693;
						shift_out14 <= X1694;
						shift_out15 <= X1695;
						i <= i + 1;
					WHEN 106 =>
						shift_out0 <= X1696;
						shift_out1 <= X1697;
						shift_out2 <= X1698;
						shift_out3 <= X1699;
						shift_out4 <= X1700;
						shift_out5 <= X1701;
						shift_out6 <= X1702;
						shift_out7 <= X1703;
						shift_out8 <= X1704;
						shift_out9 <= X1705;
						shift_out10 <= X1706;
						shift_out11 <= X1707;
						shift_out12 <= X1708;
						shift_out13 <= X1709;
						shift_out14 <= X1710;
						shift_out15 <= X1711;
						i <= i + 1;
					WHEN 107 =>
						shift_out0 <= X1712;
						shift_out1 <= X1713;
						shift_out2 <= X1714;
						shift_out3 <= X1715;
						shift_out4 <= X1716;
						shift_out5 <= X1717;
						shift_out6 <= X1718;
						shift_out7 <= X1719;
						shift_out8 <= X1720;
						shift_out9 <= X1721;
						shift_out10 <= X1722;
						shift_out11 <= X1723;
						shift_out12 <= X1724;
						shift_out13 <= X1725;
						shift_out14 <= X1726;
						shift_out15 <= X1727;
						i <= i + 1;
					WHEN 108 =>
						shift_out0 <= X1728;
						shift_out1 <= X1729;
						shift_out2 <= X1730;
						shift_out3 <= X1731;
						shift_out4 <= X1732;
						shift_out5 <= X1733;
						shift_out6 <= X1734;
						shift_out7 <= X1735;
						shift_out8 <= X1736;
						shift_out9 <= X1737;
						shift_out10 <= X1738;
						shift_out11 <= X1739;
						shift_out12 <= X1740;
						shift_out13 <= X1741;
						shift_out14 <= X1742;
						shift_out15 <= X1743;
						i <= i + 1;
					WHEN 109 =>
						shift_out0 <= X1744;
						shift_out1 <= X1745;
						shift_out2 <= X1746;
						shift_out3 <= X1747;
						shift_out4 <= X1748;
						shift_out5 <= X1749;
						shift_out6 <= X1750;
						shift_out7 <= X1751;
						shift_out8 <= X1752;
						shift_out9 <= X1753;
						shift_out10 <= X1754;
						shift_out11 <= X1755;
						shift_out12 <= X1756;
						shift_out13 <= X1757;
						shift_out14 <= X1758;
						shift_out15 <= X1759;
						i <= i + 1;
					WHEN 110 =>
						shift_out0 <= X1760;
						shift_out1 <= X1761;
						shift_out2 <= X1762;
						shift_out3 <= X1763;
						shift_out4 <= X1764;
						shift_out5 <= X1765;
						shift_out6 <= X1766;
						shift_out7 <= X1767;
						shift_out8 <= X1768;
						shift_out9 <= X1769;
						shift_out10 <= X1770;
						shift_out11 <= X1771;
						shift_out12 <= X1772;
						shift_out13 <= X1773;
						shift_out14 <= X1774;
						shift_out15 <= X1775;
						i <= i + 1;
					WHEN 111 =>
						shift_out0 <= X1776;
						shift_out1 <= X1777;
						shift_out2 <= X1778;
						shift_out3 <= X1779;
						shift_out4 <= X1780;
						shift_out5 <= X1781;
						shift_out6 <= X1782;
						shift_out7 <= X1783;
						shift_out8 <= X1784;
						shift_out9 <= X1785;
						shift_out10 <= X1786;
						shift_out11 <= X1787;
						shift_out12 <= X1788;
						shift_out13 <= X1789;
						shift_out14 <= X1790;
						shift_out15 <= X1791;
						i <= i + 1;
					WHEN 112 =>
						shift_out0 <= X1792;
						shift_out1 <= X1793;
						shift_out2 <= X1794;
						shift_out3 <= X1795;
						shift_out4 <= X1796;
						shift_out5 <= X1797;
						shift_out6 <= X1798;
						shift_out7 <= X1799;
						shift_out8 <= X1800;
						shift_out9 <= X1801;
						shift_out10 <= X1802;
						shift_out11 <= X1803;
						shift_out12 <= X1804;
						shift_out13 <= X1805;
						shift_out14 <= X1806;
						shift_out15 <= X1807;
						i <= i + 1;
					WHEN 113 =>
						shift_out0 <= X1808;
						shift_out1 <= X1809;
						shift_out2 <= X1810;
						shift_out3 <= X1811;
						shift_out4 <= X1812;
						shift_out5 <= X1813;
						shift_out6 <= X1814;
						shift_out7 <= X1815;
						shift_out8 <= X1816;
						shift_out9 <= X1817;
						shift_out10 <= X1818;
						shift_out11 <= X1819;
						shift_out12 <= X1820;
						shift_out13 <= X1821;
						shift_out14 <= X1822;
						shift_out15 <= X1823;
						i <= i + 1;
					WHEN 114 =>
						shift_out0 <= X1824;
						shift_out1 <= X1825;
						shift_out2 <= X1826;
						shift_out3 <= X1827;
						shift_out4 <= X1828;
						shift_out5 <= X1829;
						shift_out6 <= X1830;
						shift_out7 <= X1831;
						shift_out8 <= X1832;
						shift_out9 <= X1833;
						shift_out10 <= X1834;
						shift_out11 <= X1835;
						shift_out12 <= X1836;
						shift_out13 <= X1837;
						shift_out14 <= X1838;
						shift_out15 <= X1839;
						i <= i + 1;
					WHEN 115 =>
						shift_out0 <= X1840;
						shift_out1 <= X1841;
						shift_out2 <= X1842;
						shift_out3 <= X1843;
						shift_out4 <= X1844;
						shift_out5 <= X1845;
						shift_out6 <= X1846;
						shift_out7 <= X1847;
						shift_out8 <= X1848;
						shift_out9 <= X1849;
						shift_out10 <= X1850;
						shift_out11 <= X1851;
						shift_out12 <= X1852;
						shift_out13 <= X1853;
						shift_out14 <= X1854;
						shift_out15 <= X1855;
						i <= i + 1;
					WHEN 116 =>
						shift_out0 <= X1856;
						shift_out1 <= X1857;
						shift_out2 <= X1858;
						shift_out3 <= X1859;
						shift_out4 <= X1860;
						shift_out5 <= X1861;
						shift_out6 <= X1862;
						shift_out7 <= X1863;
						shift_out8 <= X1864;
						shift_out9 <= X1865;
						shift_out10 <= X1866;
						shift_out11 <= X1867;
						shift_out12 <= X1868;
						shift_out13 <= X1869;
						shift_out14 <= X1870;
						shift_out15 <= X1871;
						i <= i + 1;
					WHEN 117 =>
						shift_out0 <= X1872;
						shift_out1 <= X1873;
						shift_out2 <= X1874;
						shift_out3 <= X1875;
						shift_out4 <= X1876;
						shift_out5 <= X1877;
						shift_out6 <= X1878;
						shift_out7 <= X1879;
						shift_out8 <= X1880;
						shift_out9 <= X1881;
						shift_out10 <= X1882;
						shift_out11 <= X1883;
						shift_out12 <= X1884;
						shift_out13 <= X1885;
						shift_out14 <= X1886;
						shift_out15 <= X1887;
						i <= i + 1;
					WHEN 118 =>
						shift_out0 <= X1888;
						shift_out1 <= X1889;
						shift_out2 <= X1890;
						shift_out3 <= X1891;
						shift_out4 <= X1892;
						shift_out5 <= X1893;
						shift_out6 <= X1894;
						shift_out7 <= X1895;
						shift_out8 <= X1896;
						shift_out9 <= X1897;
						shift_out10 <= X1898;
						shift_out11 <= X1899;
						shift_out12 <= X1900;
						shift_out13 <= X1901;
						shift_out14 <= X1902;
						shift_out15 <= X1903;
						i <= i + 1;
					WHEN 119 =>
						shift_out0 <= X1904;
						shift_out1 <= X1905;
						shift_out2 <= X1906;
						shift_out3 <= X1907;
						shift_out4 <= X1908;
						shift_out5 <= X1909;
						shift_out6 <= X1910;
						shift_out7 <= X1911;
						shift_out8 <= X1912;
						shift_out9 <= X1913;
						shift_out10 <= X1914;
						shift_out11 <= X1915;
						shift_out12 <= X1916;
						shift_out13 <= X1917;
						shift_out14 <= X1918;
						shift_out15 <= X1919;
						i <= i + 1;
					WHEN 120 =>
						shift_out0 <= X1920;
						shift_out1 <= X1921;
						shift_out2 <= X1922;
						shift_out3 <= X1923;
						shift_out4 <= X1924;
						shift_out5 <= X1925;
						shift_out6 <= X1926;
						shift_out7 <= X1927;
						shift_out8 <= X1928;
						shift_out9 <= X1929;
						shift_out10 <= X1930;
						shift_out11 <= X1931;
						shift_out12 <= X1932;
						shift_out13 <= X1933;
						shift_out14 <= X1934;
						shift_out15 <= X1935;
						i <= i + 1;
					WHEN 121 =>
						shift_out0 <= X1936;
						shift_out1 <= X1937;
						shift_out2 <= X1938;
						shift_out3 <= X1939;
						shift_out4 <= X1940;
						shift_out5 <= X1941;
						shift_out6 <= X1942;
						shift_out7 <= X1943;
						shift_out8 <= X1944;
						shift_out9 <= X1945;
						shift_out10 <= X1946;
						shift_out11 <= X1947;
						shift_out12 <= X1948;
						shift_out13 <= X1949;
						shift_out14 <= X1950;
						shift_out15 <= X1951;
						i <= i + 1;
					WHEN 122 =>
						shift_out0 <= X1952;
						shift_out1 <= X1953;
						shift_out2 <= X1954;
						shift_out3 <= X1955;
						shift_out4 <= X1956;
						shift_out5 <= X1957;
						shift_out6 <= X1958;
						shift_out7 <= X1959;
						shift_out8 <= X1960;
						shift_out9 <= X1961;
						shift_out10 <= X1962;
						shift_out11 <= X1963;
						shift_out12 <= X1964;
						shift_out13 <= X1965;
						shift_out14 <= X1966;
						shift_out15 <= X1967;
						i <= i + 1;
					WHEN 123 =>
						shift_out0 <= X1968;
						shift_out1 <= X1969;
						shift_out2 <= X1970;
						shift_out3 <= X1971;
						shift_out4 <= X1972;
						shift_out5 <= X1973;
						shift_out6 <= X1974;
						shift_out7 <= X1975;
						shift_out8 <= X1976;
						shift_out9 <= X1977;
						shift_out10 <= X1978;
						shift_out11 <= X1979;
						shift_out12 <= X1980;
						shift_out13 <= X1981;
						shift_out14 <= X1982;
						shift_out15 <= X1983;
						i <= i + 1;
					WHEN 124 =>
						shift_out0 <= X1984;
						shift_out1 <= X1985;
						shift_out2 <= X1986;
						shift_out3 <= X1987;
						shift_out4 <= X1988;
						shift_out5 <= X1989;
						shift_out6 <= X1990;
						shift_out7 <= X1991;
						shift_out8 <= X1992;
						shift_out9 <= X1993;
						shift_out10 <= X1994;
						shift_out11 <= X1995;
						shift_out12 <= X1996;
						shift_out13 <= X1997;
						shift_out14 <= X1998;
						shift_out15 <= X1999;
						i <= i + 1;
					WHEN 125 =>
						shift_out0 <= X2000;
						shift_out1 <= X2001;
						shift_out2 <= X2002;
						shift_out3 <= X2003;
						shift_out4 <= X2004;
						shift_out5 <= X2005;
						shift_out6 <= X2006;
						shift_out7 <= X2007;
						shift_out8 <= X2008;
						shift_out9 <= X2009;
						shift_out10 <= X2010;
						shift_out11 <= X2011;
						shift_out12 <= X2012;
						shift_out13 <= X2013;
						shift_out14 <= X2014;
						shift_out15 <= X2015;
						i <= i + 1;
					WHEN 126 =>
						shift_out0 <= X2016;
						shift_out1 <= X2017;
						shift_out2 <= X2018;
						shift_out3 <= X2019;
						shift_out4 <= X2020;
						shift_out5 <= X2021;
						shift_out6 <= X2022;
						shift_out7 <= X2023;
						shift_out8 <= X2024;
						shift_out9 <= X2025;
						shift_out10 <= X2026;
						shift_out11 <= X2027;
						shift_out12 <= X2028;
						shift_out13 <= X2029;
						shift_out14 <= X2030;
						shift_out15 <= X2031;
						i <= i + 1;
					WHEN 127 =>
						shift_out0 <= X2032;
						shift_out1 <= X2033;
						shift_out2 <= X2034;
						shift_out3 <= X2035;
						shift_out4 <= X2036;
						shift_out5 <= X2037;
						shift_out6 <= X2038;
						shift_out7 <= X2039;
						shift_out8 <= X2040;
						shift_out9 <= X2041;
						shift_out10 <= X2042;
						shift_out11 <= X2043;
						shift_out12 <= X2044;
						shift_out13 <= X2045;
						shift_out14 <= X2046;
						shift_out15 <= X2047;
						
						i <= i + 1;	
					WHEN OTHERS =>
						reading_input <= 0;
						i <= 0;
								--do-nothing
					END CASE;
				
				WHEN OTHERS =>
				END CASE;
			END IF;
		
	END PROCESS;

END shift;
