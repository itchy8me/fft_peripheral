-- *************************************************************************
-- Author : Wernher Korff																	*
-- Function : connects the underlying architecture together and expose the *
--				FFT peripheral inputs and outputs										*
-- *************************************************************************

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

-- Top Block --
ENTITY fft_peripheral IS
	PORT(
	X0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X4 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X5 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X6 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X7 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X8 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X9 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X10 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X11 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X12 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X13 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X14 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X15 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X16 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X17 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X18 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X19 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X20 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X21 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X22 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X23 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X24 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X25 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X26 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X27 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X28 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X29 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X30 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X31 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X32 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X33 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X34 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X35 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X36 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X37 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X38 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X39 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X40 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X41 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X42 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X43 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X44 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X45 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X46 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X47 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X48 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X49 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X50 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X51 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X52 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X53 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X54 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X55 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X56 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X57 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X58 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X59 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X60 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X61 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X62 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X63 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X64 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X65 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X66 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X67 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X68 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X69 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X70 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X71 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X72 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X73 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X74 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X75 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X76 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X77 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X78 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X79 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X80 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X81 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X82 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X83 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X84 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X85 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X86 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X87 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X88 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X89 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X90 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X91 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X92 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X93 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X94 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X95 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X96 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X97 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X98 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X99 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X100 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X101 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X102 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X103 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X104 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X105 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X106 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X107 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X108 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X109 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X110 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X111 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X112 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X113 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X114 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X115 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X116 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X117 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X118 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X119 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X120 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X121 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X122 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X123 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X124 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X125 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X126 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X127 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X128 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X129 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X130 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X131 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X132 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X133 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X134 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X135 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X136 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X137 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X138 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X139 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X140 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X141 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X142 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X143 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X144 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X145 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X146 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X147 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X148 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X149 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X150 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X151 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X152 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X153 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X154 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X155 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X156 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X157 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X158 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X159 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X160 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X161 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X162 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X163 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X164 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X165 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X166 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X167 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X168 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X169 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X170 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X171 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X172 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X173 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X174 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X175 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X176 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X177 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X178 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X179 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X180 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X181 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X182 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X183 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X184 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X185 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X186 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X187 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X188 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X189 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X190 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X191 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X192 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X193 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X194 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X195 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X196 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X197 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X198 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X199 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X200 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X201 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X202 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X203 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X204 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X205 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X206 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X207 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X208 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X209 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X210 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X211 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X212 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X213 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X214 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X215 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X216 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X217 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X218 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X219 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X220 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X221 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X222 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X223 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X224 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X225 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X226 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X227 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X228 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X229 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X230 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X231 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X232 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X233 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X234 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X235 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X236 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X237 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X238 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X239 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X240 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X241 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X242 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X243 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X244 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X245 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X246 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X247 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X248 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X249 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X250 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X251 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X252 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X253 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X254 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X255 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X256 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X257 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X258 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X259 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X260 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X261 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X262 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X263 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X264 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X265 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X266 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X267 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X268 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X269 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X270 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X271 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X272 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X273 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X274 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X275 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X276 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X277 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X278 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X279 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X280 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X281 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X282 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X283 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X284 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X285 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X286 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X287 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X288 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X289 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X290 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X291 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X292 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X293 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X294 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X295 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X296 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X297 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X298 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X299 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X300 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X301 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X302 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X303 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X304 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X305 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X306 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X307 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X308 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X309 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X310 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X311 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X312 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X313 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X314 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X315 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X316 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X317 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X318 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X319 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X320 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X321 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X322 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X323 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X324 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X325 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X326 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X327 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X328 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X329 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X330 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X331 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X332 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X333 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X334 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X335 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X336 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X337 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X338 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X339 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X340 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X341 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X342 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X343 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X344 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X345 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X346 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X347 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X348 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X349 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X350 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X351 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X352 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X353 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X354 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X355 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X356 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X357 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X358 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X359 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X360 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X361 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X362 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X363 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X364 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X365 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X366 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X367 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X368 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X369 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X370 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X371 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X372 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X373 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X374 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X375 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X376 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X377 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X378 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X379 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X380 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X381 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X382 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X383 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X384 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X385 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X386 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X387 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X388 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X389 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X390 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X391 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X392 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X393 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X394 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X395 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X396 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X397 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X398 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X399 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X400 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X401 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X402 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X403 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X404 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X405 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X406 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X407 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X408 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X409 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X410 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X411 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X412 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X413 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X414 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X415 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X416 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X417 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X418 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X419 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X420 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X421 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X422 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X423 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X424 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X425 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X426 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X427 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X428 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X429 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X430 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X431 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X432 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X433 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X434 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X435 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X436 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X437 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X438 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X439 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X440 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X441 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X442 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X443 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X444 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X445 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X446 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X447 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X448 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X449 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X450 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X451 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X452 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X453 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X454 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X455 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X456 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X457 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X458 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X459 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X460 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X461 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X462 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X463 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X464 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X465 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X466 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X467 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X468 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X469 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X470 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X471 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X472 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X473 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X474 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X475 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X476 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X477 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X478 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X479 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X480 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X481 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X482 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X483 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X484 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X485 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X486 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X487 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X488 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X489 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X490 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X491 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X492 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X493 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X494 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X495 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X496 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X497 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X498 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X499 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X500 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X501 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X502 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X503 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X504 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X505 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X506 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X507 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X508 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X509 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X510 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X511 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X512 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X513 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X514 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X515 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X516 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X517 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X518 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X519 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X520 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X521 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X522 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X523 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X524 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X525 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X526 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X527 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X528 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X529 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X530 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X531 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X532 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X533 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X534 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X535 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X536 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X537 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X538 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X539 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X540 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X541 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X542 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X543 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X544 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X545 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X546 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X547 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X548 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X549 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X550 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X551 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X552 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X553 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X554 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X555 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X556 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X557 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X558 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X559 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X560 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X561 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X562 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X563 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X564 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X565 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X566 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X567 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X568 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X569 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X570 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X571 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X572 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X573 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X574 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X575 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X576 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X577 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X578 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X579 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X580 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X581 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X582 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X583 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X584 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X585 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X586 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X587 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X588 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X589 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X590 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X591 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X592 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X593 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X594 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X595 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X596 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X597 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X598 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X599 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X600 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X601 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X602 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X603 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X604 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X605 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X606 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X607 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X608 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X609 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X610 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X611 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X612 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X613 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X614 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X615 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X616 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X617 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X618 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X619 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X620 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X621 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X622 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X623 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X624 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X625 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X626 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X627 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X628 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X629 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X630 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X631 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X632 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X633 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X634 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X635 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X636 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X637 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X638 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X639 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X640 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X641 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X642 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X643 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X644 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X645 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X646 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X647 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X648 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X649 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X650 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X651 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X652 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X653 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X654 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X655 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X656 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X657 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X658 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X659 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X660 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X661 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X662 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X663 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X664 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X665 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X666 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X667 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X668 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X669 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X670 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X671 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X672 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X673 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X674 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X675 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X676 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X677 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X678 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X679 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X680 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X681 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X682 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X683 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X684 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X685 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X686 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X687 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X688 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X689 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X690 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X691 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X692 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X693 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X694 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X695 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X696 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X697 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X698 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X699 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X700 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X701 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X702 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X703 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X704 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X705 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X706 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X707 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X708 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X709 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X710 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X711 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X712 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X713 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X714 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X715 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X716 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X717 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X718 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X719 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X720 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X721 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X722 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X723 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X724 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X725 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X726 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X727 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X728 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X729 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X730 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X731 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X732 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X733 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X734 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X735 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X736 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X737 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X738 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X739 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X740 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X741 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X742 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X743 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X744 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X745 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X746 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X747 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X748 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X749 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X750 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X751 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X752 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X753 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X754 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X755 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X756 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X757 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X758 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X759 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X760 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X761 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X762 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X763 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X764 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X765 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X766 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X767 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X768 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X769 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X770 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X771 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X772 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X773 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X774 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X775 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X776 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X777 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X778 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X779 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X780 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X781 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X782 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X783 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X784 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X785 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X786 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X787 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X788 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X789 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X790 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X791 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X792 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X793 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X794 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X795 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X796 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X797 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X798 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X799 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X800 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X801 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X802 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X803 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X804 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X805 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X806 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X807 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X808 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X809 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X810 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X811 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X812 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X813 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X814 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X815 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X816 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X817 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X818 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X819 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X820 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X821 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X822 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X823 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X824 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X825 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X826 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X827 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X828 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X829 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X830 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X831 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X832 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X833 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X834 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X835 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X836 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X837 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X838 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X839 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X840 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X841 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X842 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X843 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X844 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X845 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X846 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X847 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X848 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X849 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X850 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X851 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X852 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X853 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X854 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X855 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X856 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X857 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X858 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X859 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X860 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X861 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X862 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X863 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X864 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X865 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X866 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X867 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X868 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X869 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X870 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X871 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X872 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X873 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X874 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X875 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X876 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X877 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X878 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X879 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X880 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X881 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X882 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X883 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X884 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X885 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X886 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X887 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X888 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X889 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X890 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X891 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X892 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X893 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X894 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X895 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X896 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X897 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X898 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X899 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X900 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X901 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X902 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X903 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X904 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X905 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X906 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X907 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X908 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X909 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X910 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X911 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X912 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X913 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X914 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X915 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X916 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X917 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X918 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X919 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X920 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X921 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X922 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X923 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X924 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X925 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X926 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X927 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X928 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X929 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X930 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X931 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X932 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X933 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X934 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X935 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X936 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X937 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X938 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X939 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X940 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X941 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X942 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X943 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X944 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X945 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X946 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X947 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X948 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X949 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X950 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X951 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X952 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X953 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X954 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X955 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X956 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X957 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X958 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X959 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X960 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X961 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X962 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X963 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X964 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X965 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X966 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X967 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X968 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X969 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X970 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X971 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X972 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X973 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X974 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X975 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X976 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X977 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X978 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X979 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X980 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X981 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X982 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X983 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X984 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X985 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X986 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X987 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X988 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X989 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X990 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X991 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X992 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X993 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X994 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X995 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X996 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X997 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X998 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X999 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1000 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1001 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1002 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1003 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1004 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1005 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1006 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1007 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1008 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1009 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1010 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1011 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1012 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1013 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1014 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1015 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1016 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1017 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1018 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1019 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1020 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1021 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1022 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1023 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1024 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1025 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1026 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1027 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1028 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1029 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1030 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1031 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1032 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1033 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1034 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1035 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1036 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1037 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1038 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1039 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1040 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1041 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1042 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1043 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1044 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1045 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1046 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1047 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1048 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1049 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1050 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1051 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1052 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1053 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1054 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1055 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1056 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1057 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1058 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1059 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1060 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1061 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1062 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1063 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1064 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1065 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1066 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1067 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1068 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1069 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1070 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1071 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1072 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1073 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1074 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1075 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1076 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1077 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1078 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1079 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1080 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1081 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1082 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1083 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1084 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1085 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1086 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1087 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1088 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1089 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1090 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1091 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1092 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1093 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1094 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1095 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1096 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1097 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1098 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1099 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1100 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1101 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1102 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1103 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1104 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1105 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1106 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1107 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1108 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1109 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1110 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1111 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1112 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1113 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1114 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1115 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1116 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1117 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1118 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1119 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1120 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1121 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1122 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1123 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1124 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1125 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1126 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1127 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1128 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1129 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1130 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1131 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1132 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1133 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1134 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1135 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1136 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1137 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1138 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1139 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1140 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1141 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1142 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1143 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1144 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1145 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1146 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1147 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1148 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1149 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1150 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1151 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1152 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1153 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1154 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1155 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1156 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1157 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1158 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1159 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1160 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1161 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1162 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1163 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1164 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1165 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1166 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1167 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1168 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1169 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1170 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1171 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1172 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1173 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1174 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1175 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1176 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1177 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1178 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1179 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1180 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1181 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1182 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1183 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1184 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1185 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1186 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1187 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1188 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1189 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1190 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1191 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1192 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1193 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1194 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1195 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1196 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1197 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1198 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1199 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1200 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1201 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1202 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1203 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1204 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1205 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1206 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1207 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1208 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1209 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1210 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1211 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1212 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1213 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1214 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1215 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1216 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1217 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1218 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1219 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1220 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1221 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1222 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1223 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1224 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1225 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1226 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1227 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1228 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1229 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1230 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1231 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1232 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1233 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1234 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1235 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1236 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1237 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1238 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1239 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1240 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1241 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1242 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1243 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1244 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1245 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1246 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1247 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1248 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1249 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1250 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1251 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1252 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1253 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1254 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1255 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1256 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1257 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1258 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1259 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1260 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1261 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1262 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1263 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1264 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1265 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1266 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1267 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1268 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1269 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1270 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1271 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1272 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1273 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1274 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1275 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1276 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1277 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1278 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1279 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1280 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1281 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1282 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1283 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1284 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1285 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1286 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1287 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1288 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1289 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1290 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1291 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1292 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1293 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1294 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1295 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1296 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1297 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1298 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1299 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1300 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1301 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1302 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1303 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1304 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1305 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1306 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1307 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1308 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1309 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1310 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1311 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1312 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1313 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1314 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1315 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1316 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1317 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1318 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1319 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1320 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1321 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1322 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1323 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1324 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1325 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1326 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1327 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1328 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1329 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1330 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1331 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1332 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1333 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1334 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1335 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1336 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1337 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1338 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1339 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1340 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1341 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1342 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1343 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1344 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1345 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1346 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1347 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1348 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1349 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1350 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1351 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1352 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1353 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1354 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1355 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1356 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1357 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1358 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1359 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1360 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1361 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1362 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1363 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1364 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1365 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1366 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1367 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1368 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1369 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1370 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1371 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1372 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1373 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1374 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1375 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1376 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1377 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1378 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1379 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1380 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1381 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1382 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1383 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1384 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1385 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1386 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1387 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1388 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1389 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1390 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1391 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1392 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1393 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1394 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1395 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1396 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1397 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1398 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1399 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1400 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1401 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1402 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1403 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1404 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1405 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1406 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1407 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1408 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1409 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1410 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1411 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1412 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1413 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1414 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1415 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1416 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1417 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1418 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1419 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1420 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1421 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1422 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1423 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1424 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1425 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1426 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1427 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1428 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1429 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1430 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1431 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1432 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1433 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1434 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1435 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1436 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1437 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1438 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1439 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1440 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1441 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1442 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1443 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1444 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1445 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1446 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1447 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1448 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1449 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1450 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1451 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1452 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1453 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1454 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1455 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1456 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1457 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1458 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1459 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1460 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1461 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1462 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1463 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1464 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1465 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1466 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1467 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1468 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1469 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1470 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1471 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1472 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1473 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1474 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1475 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1476 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1477 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1478 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1479 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1480 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1481 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1482 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1483 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1484 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1485 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1486 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1487 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1488 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1489 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1490 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1491 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1492 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1493 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1494 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1495 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1496 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1497 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1498 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1499 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1500 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1501 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1502 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1503 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1504 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1505 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1506 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1507 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1508 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1509 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1510 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1511 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1512 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1513 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1514 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1515 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1516 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1517 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1518 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1519 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1520 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1521 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1522 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1523 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1524 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1525 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1526 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1527 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1528 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1529 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1530 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1531 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1532 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1533 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1534 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1535 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1536 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1537 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1538 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1539 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1540 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1541 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1542 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1543 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1544 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1545 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1546 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1547 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1548 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1549 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1550 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1551 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1552 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1553 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1554 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1555 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1556 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1557 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1558 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1559 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1560 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1561 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1562 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1563 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1564 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1565 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1566 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1567 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1568 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1569 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1570 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1571 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1572 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1573 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1574 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1575 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1576 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1577 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1578 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1579 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1580 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1581 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1582 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1583 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1584 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1585 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1586 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1587 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1588 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1589 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1590 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1591 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1592 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1593 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1594 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1595 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1596 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1597 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1598 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1599 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1600 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1601 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1602 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1603 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1604 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1605 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1606 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1607 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1608 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1609 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1610 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1611 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1612 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1613 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1614 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1615 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1616 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1617 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1618 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1619 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1620 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1621 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1622 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1623 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1624 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1625 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1626 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1627 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1628 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1629 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1630 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1631 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1632 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1633 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1634 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1635 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1636 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1637 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1638 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1639 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1640 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1641 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1642 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1643 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1644 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1645 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1646 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1647 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1648 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1649 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1650 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1651 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1652 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1653 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1654 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1655 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1656 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1657 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1658 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1659 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1660 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1661 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1662 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1663 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1664 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1665 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1666 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1667 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1668 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1669 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1670 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1671 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1672 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1673 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1674 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1675 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1676 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1677 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1678 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1679 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1680 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1681 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1682 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1683 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1684 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1685 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1686 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1687 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1688 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1689 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1690 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1691 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1692 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1693 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1694 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1695 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1696 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1697 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1698 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1699 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1700 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1701 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1702 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1703 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1704 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1705 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1706 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1707 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1708 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1709 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1710 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1711 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1712 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1713 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1714 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1715 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1716 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1717 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1718 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1719 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1720 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1721 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1722 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1723 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1724 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1725 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1726 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1727 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1728 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1729 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1730 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1731 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1732 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1733 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1734 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1735 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1736 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1737 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1738 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1739 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1740 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1741 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1742 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1743 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1744 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1745 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1746 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1747 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1748 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1749 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1750 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1751 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1752 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1753 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1754 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1755 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1756 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1757 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1758 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1759 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1760 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1761 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1762 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1763 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1764 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1765 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1766 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1767 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1768 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1769 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1770 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1771 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1772 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1773 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1774 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1775 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1776 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1777 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1778 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1779 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1780 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1781 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1782 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1783 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1784 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1785 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1786 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1787 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1788 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1789 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1790 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1791 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1792 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1793 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1794 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1795 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1796 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1797 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1798 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1799 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1800 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1801 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1802 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1803 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1804 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1805 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1806 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1807 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1808 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1809 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1810 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1811 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1812 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1813 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1814 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1815 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1816 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1817 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1818 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1819 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1820 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1821 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1822 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1823 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1824 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1825 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1826 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1827 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1828 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1829 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1830 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1831 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1832 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1833 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1834 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1835 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1836 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1837 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1838 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1839 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1840 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1841 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1842 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1843 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1844 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1845 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1846 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1847 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1848 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1849 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1850 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1851 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1852 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1853 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1854 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1855 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1856 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1857 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1858 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1859 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1860 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1861 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1862 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1863 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1864 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1865 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1866 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1867 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1868 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1869 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1870 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1871 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1872 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1873 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1874 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1875 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1876 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1877 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1878 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1879 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1880 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1881 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1882 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1883 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1884 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1885 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1886 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1887 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1888 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1889 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1890 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1891 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1892 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1893 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1894 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1895 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1896 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1897 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1898 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1899 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1900 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1901 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1902 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1903 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1904 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1905 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1906 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1907 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1908 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1909 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1910 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1911 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1912 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1913 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1914 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1915 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1916 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1917 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1918 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1919 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1920 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1921 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1922 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1923 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1924 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1925 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1926 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1927 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1928 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1929 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1930 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1931 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1932 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1933 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1934 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1935 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1936 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1937 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1938 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1939 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1940 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1941 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1942 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1943 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1944 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1945 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1946 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1947 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1948 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1949 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1950 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1951 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1952 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1953 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1954 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1955 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1956 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1957 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1958 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1959 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1960 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1961 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1962 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1963 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1964 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1965 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1966 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1967 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1968 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1969 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1970 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1971 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1972 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1973 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1974 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1975 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1976 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1977 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1978 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1979 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1980 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1981 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1982 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1983 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1984 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1985 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1986 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1987 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1988 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1989 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1990 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1991 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1992 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1993 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1994 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1995 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1996 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1997 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1998 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X1999 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2000 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2001 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2002 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2003 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2004 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2005 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2006 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2007 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2008 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2009 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2010 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2011 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2012 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2013 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2014 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2015 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2016 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2017 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2018 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2019 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2020 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2021 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2022 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2023 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2024 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2025 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2026 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2027 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2028 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2029 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2030 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2031 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2032 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2033 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2034 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2035 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2036 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2037 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2038 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2039 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2040 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2041 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2042 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2043 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2044 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2045 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2046 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	X2047 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	
	samples_ready : IN STD_LOGIC := '0';	-- sampler has 2048 samples ready
	clk : IN STD_LOGIC := '0';
	fft_finished : OUT STD_LOGIC := '0';	-- the system is idle / can receive data
	
	busy : IN STD_LOGIC := '0';	-- receiving side status
	data_ready : OUT STD_LOGIC := '0'; -- the FFT has data ready for output / cycle data
	
	-- data ouput for interfacing device 64 sets of 16 
	V0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	V1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	V2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	V3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	V4 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	V5 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	V6 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	V7 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	V8 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	V9 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	V10 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	V11 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	V12 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	V13 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	V14 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	V15 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000");
END fft_peripheral;


-- mapping together of components --
ARCHITECTURE interconnect OF fft_peripheral IS
	
	-- the fft block --
	COMPONENT dft_top
	PORT (
		clk : IN STD_LOGIC := '0';
		reset : IN STD_LOGIC := '0';
		next_in : IN STD_LOGIC := '0';
		next_out : OUT STD_LOGIC := '0';
		X0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X4 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X5 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X6 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X7 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X8 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X9 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X10 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X11 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X12 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X13 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X14 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X15 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X16 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X17 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X18 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X19 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X20 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X21 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X22 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X23 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X24 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X25 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X26 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X27 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X28 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X29 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X30 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X31 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		
		Y0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y4 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y5 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y6 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y7 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y8 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y9 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y10 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y11 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y12 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y13 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y14 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y15 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y16 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y17 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y18 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y19 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y20 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y21 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y22 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y23 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y24 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y25 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y26 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y27 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y28 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y29 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y30 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		Y31 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000");
	END COMPONENT; -- dft_top
	
	-- controls the clock to th efft and input shifter, when busy is '0' and converting '0' then clock is active,
	-- otherwise it is inactive
	COMPONENT clock_control
	PORT(
		disable_1 : IN STD_LOGIC := '0';
		disable_2: IN STD_LOGIC := '0';
		clock : IN STD_LOGIC := '0';
		
		controlled_clock : OUT STD_LOGIC := '0');
	END COMPONENT; -- clock_control
	
	
	-- divvides 2048 samples into 64 sets of 16 samples each --
	COMPONENT c_2048to16x128_shifter
		PORT (
		X0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X4 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X5 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X6 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X7 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X8 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X9 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X10 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X11 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X12 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X13 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X14 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X15 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X16 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X17 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X18 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X19 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X20 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X21 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X22 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X23 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X24 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X25 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X26 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X27 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X28 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X29 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X30 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X31 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X32 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X33 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X34 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X35 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X36 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X37 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X38 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X39 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X40 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X41 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X42 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X43 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X44 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X45 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X46 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X47 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X48 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X49 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X50 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X51 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X52 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X53 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X54 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X55 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X56 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X57 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X58 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X59 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X60 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X61 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X62 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X63 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X64 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X65 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X66 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X67 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X68 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X69 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X70 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X71 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X72 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X73 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X74 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X75 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X76 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X77 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X78 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X79 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X80 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X81 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X82 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X83 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X84 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X85 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X86 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X87 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X88 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X89 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X90 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X91 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X92 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X93 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X94 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X95 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X96 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X97 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X98 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X99 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X100 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X101 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X102 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X103 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X104 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X105 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X106 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X107 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X108 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X109 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X110 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X111 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X112 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X113 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X114 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X115 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X116 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X117 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X118 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X119 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X120 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X121 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X122 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X123 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X124 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X125 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X126 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X127 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X128 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X129 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X130 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X131 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X132 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X133 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X134 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X135 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X136 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X137 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X138 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X139 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X140 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X141 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X142 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X143 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X144 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X145 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X146 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X147 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X148 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X149 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X150 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X151 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X152 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X153 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X154 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X155 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X156 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X157 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X158 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X159 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X160 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X161 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X162 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X163 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X164 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X165 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X166 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X167 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X168 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X169 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X170 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X171 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X172 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X173 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X174 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X175 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X176 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X177 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X178 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X179 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X180 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X181 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X182 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X183 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X184 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X185 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X186 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X187 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X188 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X189 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X190 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X191 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X192 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X193 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X194 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X195 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X196 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X197 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X198 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X199 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X200 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X201 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X202 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X203 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X204 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X205 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X206 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X207 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X208 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X209 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X210 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X211 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X212 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X213 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X214 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X215 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X216 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X217 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X218 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X219 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X220 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X221 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X222 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X223 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X224 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X225 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X226 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X227 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X228 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X229 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X230 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X231 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X232 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X233 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X234 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X235 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X236 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X237 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X238 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X239 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X240 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X241 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X242 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X243 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X244 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X245 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X246 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X247 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X248 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X249 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X250 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X251 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X252 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X253 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X254 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X255 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X256 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X257 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X258 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X259 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X260 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X261 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X262 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X263 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X264 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X265 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X266 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X267 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X268 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X269 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X270 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X271 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X272 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X273 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X274 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X275 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X276 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X277 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X278 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X279 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X280 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X281 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X282 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X283 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X284 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X285 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X286 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X287 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X288 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X289 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X290 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X291 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X292 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X293 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X294 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X295 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X296 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X297 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X298 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X299 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X300 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X301 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X302 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X303 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X304 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X305 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X306 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X307 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X308 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X309 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X310 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X311 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X312 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X313 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X314 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X315 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X316 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X317 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X318 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X319 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X320 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X321 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X322 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X323 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X324 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X325 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X326 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X327 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X328 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X329 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X330 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X331 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X332 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X333 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X334 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X335 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X336 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X337 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X338 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X339 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X340 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X341 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X342 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X343 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X344 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X345 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X346 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X347 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X348 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X349 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X350 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X351 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X352 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X353 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X354 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X355 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X356 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X357 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X358 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X359 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X360 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X361 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X362 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X363 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X364 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X365 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X366 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X367 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X368 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X369 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X370 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X371 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X372 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X373 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X374 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X375 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X376 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X377 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X378 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X379 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X380 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X381 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X382 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X383 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X384 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X385 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X386 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X387 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X388 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X389 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X390 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X391 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X392 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X393 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X394 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X395 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X396 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X397 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X398 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X399 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X400 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X401 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X402 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X403 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X404 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X405 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X406 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X407 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X408 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X409 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X410 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X411 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X412 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X413 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X414 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X415 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X416 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X417 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X418 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X419 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X420 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X421 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X422 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X423 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X424 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X425 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X426 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X427 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X428 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X429 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X430 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X431 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X432 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X433 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X434 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X435 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X436 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X437 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X438 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X439 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X440 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X441 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X442 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X443 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X444 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X445 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X446 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X447 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X448 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X449 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X450 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X451 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X452 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X453 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X454 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X455 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X456 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X457 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X458 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X459 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X460 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X461 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X462 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X463 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X464 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X465 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X466 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X467 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X468 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X469 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X470 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X471 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X472 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X473 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X474 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X475 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X476 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X477 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X478 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X479 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X480 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X481 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X482 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X483 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X484 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X485 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X486 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X487 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X488 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X489 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X490 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X491 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X492 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X493 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X494 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X495 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X496 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X497 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X498 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X499 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X500 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X501 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X502 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X503 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X504 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X505 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X506 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X507 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X508 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X509 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X510 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X511 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X512 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X513 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X514 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X515 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X516 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X517 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X518 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X519 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X520 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X521 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X522 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X523 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X524 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X525 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X526 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X527 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X528 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X529 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X530 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X531 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X532 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X533 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X534 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X535 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X536 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X537 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X538 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X539 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X540 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X541 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X542 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X543 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X544 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X545 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X546 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X547 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X548 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X549 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X550 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X551 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X552 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X553 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X554 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X555 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X556 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X557 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X558 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X559 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X560 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X561 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X562 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X563 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X564 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X565 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X566 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X567 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X568 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X569 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X570 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X571 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X572 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X573 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X574 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X575 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X576 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X577 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X578 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X579 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X580 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X581 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X582 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X583 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X584 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X585 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X586 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X587 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X588 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X589 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X590 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X591 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X592 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X593 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X594 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X595 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X596 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X597 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X598 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X599 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X600 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X601 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X602 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X603 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X604 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X605 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X606 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X607 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X608 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X609 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X610 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X611 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X612 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X613 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X614 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X615 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X616 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X617 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X618 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X619 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X620 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X621 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X622 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X623 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X624 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X625 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X626 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X627 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X628 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X629 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X630 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X631 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X632 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X633 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X634 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X635 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X636 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X637 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X638 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X639 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X640 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X641 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X642 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X643 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X644 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X645 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X646 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X647 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X648 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X649 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X650 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X651 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X652 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X653 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X654 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X655 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X656 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X657 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X658 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X659 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X660 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X661 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X662 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X663 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X664 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X665 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X666 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X667 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X668 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X669 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X670 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X671 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X672 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X673 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X674 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X675 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X676 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X677 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X678 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X679 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X680 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X681 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X682 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X683 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X684 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X685 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X686 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X687 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X688 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X689 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X690 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X691 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X692 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X693 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X694 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X695 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X696 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X697 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X698 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X699 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X700 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X701 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X702 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X703 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X704 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X705 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X706 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X707 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X708 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X709 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X710 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X711 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X712 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X713 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X714 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X715 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X716 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X717 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X718 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X719 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X720 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X721 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X722 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X723 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X724 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X725 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X726 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X727 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X728 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X729 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X730 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X731 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X732 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X733 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X734 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X735 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X736 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X737 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X738 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X739 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X740 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X741 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X742 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X743 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X744 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X745 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X746 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X747 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X748 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X749 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X750 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X751 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X752 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X753 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X754 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X755 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X756 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X757 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X758 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X759 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X760 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X761 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X762 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X763 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X764 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X765 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X766 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X767 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X768 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X769 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X770 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X771 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X772 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X773 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X774 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X775 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X776 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X777 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X778 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X779 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X780 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X781 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X782 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X783 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X784 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X785 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X786 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X787 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X788 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X789 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X790 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X791 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X792 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X793 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X794 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X795 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X796 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X797 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X798 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X799 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X800 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X801 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X802 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X803 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X804 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X805 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X806 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X807 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X808 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X809 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X810 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X811 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X812 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X813 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X814 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X815 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X816 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X817 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X818 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X819 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X820 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X821 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X822 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X823 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X824 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X825 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X826 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X827 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X828 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X829 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X830 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X831 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X832 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X833 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X834 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X835 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X836 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X837 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X838 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X839 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X840 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X841 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X842 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X843 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X844 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X845 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X846 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X847 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X848 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X849 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X850 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X851 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X852 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X853 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X854 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X855 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X856 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X857 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X858 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X859 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X860 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X861 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X862 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X863 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X864 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X865 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X866 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X867 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X868 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X869 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X870 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X871 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X872 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X873 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X874 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X875 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X876 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X877 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X878 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X879 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X880 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X881 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X882 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X883 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X884 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X885 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X886 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X887 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X888 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X889 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X890 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X891 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X892 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X893 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X894 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X895 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X896 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X897 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X898 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X899 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X900 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X901 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X902 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X903 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X904 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X905 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X906 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X907 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X908 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X909 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X910 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X911 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X912 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X913 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X914 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X915 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X916 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X917 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X918 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X919 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X920 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X921 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X922 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X923 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X924 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X925 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X926 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X927 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X928 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X929 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X930 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X931 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X932 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X933 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X934 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X935 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X936 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X937 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X938 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X939 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X940 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X941 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X942 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X943 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X944 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X945 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X946 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X947 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X948 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X949 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X950 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X951 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X952 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X953 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X954 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X955 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X956 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X957 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X958 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X959 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X960 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X961 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X962 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X963 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X964 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X965 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X966 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X967 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X968 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X969 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X970 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X971 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X972 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X973 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X974 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X975 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X976 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X977 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X978 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X979 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X980 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X981 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X982 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X983 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X984 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X985 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X986 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X987 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X988 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X989 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X990 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X991 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X992 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X993 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X994 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X995 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X996 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X997 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X998 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X999 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1000 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1001 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1002 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1003 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1004 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1005 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1006 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1007 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1008 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1009 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1010 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1011 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1012 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1013 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1014 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1015 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1016 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1017 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1018 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1019 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1020 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1021 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1022 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1023 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1024 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1025 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1026 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1027 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1028 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1029 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1030 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1031 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1032 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1033 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1034 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1035 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1036 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1037 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1038 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1039 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1040 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1041 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1042 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1043 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1044 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1045 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1046 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1047 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1048 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1049 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1050 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1051 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1052 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1053 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1054 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1055 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1056 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1057 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1058 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1059 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1060 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1061 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1062 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1063 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1064 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1065 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1066 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1067 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1068 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1069 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1070 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1071 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1072 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1073 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1074 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1075 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1076 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1077 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1078 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1079 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1080 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1081 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1082 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1083 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1084 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1085 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1086 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1087 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1088 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1089 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1090 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1091 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1092 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1093 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1094 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1095 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1096 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1097 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1098 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1099 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1100 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1101 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1102 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1103 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1104 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1105 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1106 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1107 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1108 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1109 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1110 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1111 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1112 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1113 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1114 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1115 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1116 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1117 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1118 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1119 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1120 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1121 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1122 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1123 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1124 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1125 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1126 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1127 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1128 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1129 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1130 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1131 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1132 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1133 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1134 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1135 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1136 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1137 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1138 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1139 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1140 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1141 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1142 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1143 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1144 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1145 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1146 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1147 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1148 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1149 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1150 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1151 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1152 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1153 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1154 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1155 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1156 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1157 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1158 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1159 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1160 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1161 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1162 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1163 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1164 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1165 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1166 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1167 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1168 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1169 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1170 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1171 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1172 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1173 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1174 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1175 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1176 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1177 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1178 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1179 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1180 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1181 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1182 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1183 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1184 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1185 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1186 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1187 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1188 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1189 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1190 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1191 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1192 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1193 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1194 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1195 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1196 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1197 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1198 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1199 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1200 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1201 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1202 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1203 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1204 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1205 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1206 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1207 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1208 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1209 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1210 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1211 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1212 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1213 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1214 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1215 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1216 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1217 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1218 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1219 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1220 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1221 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1222 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1223 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1224 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1225 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1226 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1227 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1228 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1229 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1230 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1231 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1232 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1233 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1234 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1235 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1236 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1237 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1238 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1239 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1240 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1241 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1242 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1243 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1244 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1245 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1246 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1247 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1248 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1249 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1250 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1251 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1252 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1253 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1254 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1255 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1256 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1257 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1258 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1259 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1260 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1261 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1262 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1263 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1264 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1265 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1266 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1267 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1268 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1269 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1270 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1271 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1272 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1273 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1274 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1275 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1276 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1277 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1278 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1279 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1280 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1281 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1282 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1283 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1284 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1285 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1286 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1287 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1288 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1289 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1290 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1291 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1292 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1293 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1294 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1295 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1296 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1297 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1298 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1299 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1300 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1301 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1302 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1303 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1304 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1305 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1306 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1307 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1308 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1309 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1310 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1311 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1312 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1313 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1314 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1315 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1316 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1317 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1318 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1319 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1320 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1321 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1322 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1323 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1324 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1325 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1326 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1327 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1328 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1329 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1330 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1331 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1332 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1333 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1334 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1335 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1336 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1337 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1338 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1339 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1340 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1341 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1342 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1343 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1344 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1345 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1346 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1347 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1348 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1349 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1350 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1351 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1352 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1353 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1354 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1355 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1356 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1357 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1358 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1359 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1360 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1361 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1362 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1363 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1364 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1365 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1366 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1367 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1368 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1369 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1370 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1371 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1372 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1373 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1374 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1375 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1376 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1377 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1378 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1379 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1380 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1381 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1382 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1383 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1384 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1385 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1386 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1387 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1388 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1389 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1390 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1391 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1392 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1393 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1394 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1395 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1396 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1397 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1398 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1399 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1400 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1401 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1402 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1403 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1404 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1405 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1406 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1407 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1408 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1409 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1410 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1411 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1412 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1413 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1414 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1415 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1416 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1417 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1418 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1419 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1420 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1421 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1422 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1423 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1424 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1425 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1426 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1427 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1428 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1429 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1430 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1431 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1432 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1433 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1434 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1435 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1436 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1437 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1438 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1439 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1440 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1441 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1442 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1443 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1444 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1445 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1446 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1447 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1448 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1449 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1450 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1451 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1452 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1453 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1454 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1455 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1456 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1457 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1458 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1459 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1460 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1461 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1462 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1463 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1464 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1465 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1466 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1467 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1468 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1469 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1470 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1471 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1472 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1473 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1474 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1475 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1476 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1477 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1478 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1479 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1480 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1481 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1482 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1483 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1484 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1485 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1486 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1487 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1488 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1489 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1490 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1491 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1492 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1493 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1494 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1495 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1496 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1497 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1498 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1499 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1500 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1501 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1502 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1503 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1504 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1505 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1506 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1507 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1508 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1509 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1510 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1511 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1512 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1513 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1514 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1515 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1516 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1517 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1518 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1519 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1520 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1521 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1522 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1523 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1524 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1525 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1526 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1527 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1528 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1529 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1530 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1531 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1532 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1533 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1534 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1535 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1536 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1537 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1538 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1539 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1540 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1541 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1542 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1543 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1544 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1545 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1546 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1547 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1548 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1549 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1550 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1551 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1552 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1553 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1554 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1555 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1556 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1557 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1558 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1559 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1560 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1561 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1562 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1563 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1564 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1565 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1566 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1567 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1568 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1569 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1570 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1571 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1572 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1573 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1574 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1575 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1576 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1577 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1578 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1579 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1580 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1581 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1582 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1583 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1584 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1585 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1586 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1587 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1588 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1589 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1590 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1591 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1592 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1593 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1594 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1595 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1596 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1597 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1598 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1599 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1600 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1601 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1602 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1603 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1604 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1605 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1606 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1607 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1608 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1609 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1610 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1611 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1612 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1613 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1614 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1615 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1616 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1617 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1618 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1619 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1620 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1621 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1622 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1623 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1624 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1625 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1626 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1627 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1628 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1629 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1630 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1631 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1632 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1633 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1634 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1635 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1636 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1637 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1638 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1639 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1640 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1641 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1642 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1643 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1644 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1645 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1646 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1647 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1648 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1649 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1650 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1651 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1652 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1653 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1654 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1655 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1656 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1657 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1658 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1659 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1660 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1661 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1662 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1663 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1664 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1665 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1666 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1667 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1668 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1669 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1670 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1671 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1672 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1673 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1674 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1675 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1676 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1677 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1678 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1679 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1680 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1681 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1682 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1683 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1684 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1685 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1686 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1687 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1688 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1689 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1690 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1691 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1692 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1693 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1694 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1695 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1696 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1697 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1698 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1699 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1700 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1701 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1702 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1703 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1704 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1705 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1706 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1707 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1708 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1709 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1710 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1711 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1712 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1713 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1714 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1715 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1716 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1717 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1718 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1719 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1720 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1721 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1722 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1723 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1724 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1725 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1726 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1727 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1728 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1729 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1730 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1731 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1732 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1733 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1734 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1735 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1736 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1737 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1738 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1739 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1740 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1741 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1742 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1743 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1744 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1745 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1746 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1747 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1748 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1749 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1750 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1751 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1752 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1753 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1754 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1755 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1756 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1757 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1758 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1759 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1760 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1761 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1762 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1763 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1764 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1765 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1766 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1767 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1768 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1769 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1770 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1771 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1772 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1773 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1774 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1775 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1776 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1777 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1778 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1779 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1780 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1781 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1782 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1783 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1784 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1785 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1786 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1787 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1788 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1789 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1790 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1791 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1792 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1793 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1794 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1795 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1796 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1797 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1798 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1799 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1800 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1801 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1802 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1803 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1804 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1805 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1806 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1807 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1808 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1809 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1810 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1811 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1812 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1813 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1814 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1815 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1816 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1817 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1818 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1819 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1820 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1821 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1822 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1823 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1824 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1825 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1826 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1827 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1828 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1829 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1830 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1831 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1832 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1833 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1834 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1835 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1836 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1837 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1838 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1839 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1840 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1841 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1842 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1843 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1844 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1845 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1846 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1847 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1848 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1849 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1850 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1851 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1852 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1853 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1854 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1855 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1856 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1857 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1858 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1859 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1860 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1861 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1862 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1863 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1864 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1865 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1866 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1867 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1868 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1869 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1870 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1871 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1872 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1873 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1874 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1875 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1876 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1877 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1878 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1879 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1880 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1881 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1882 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1883 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1884 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1885 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1886 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1887 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1888 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1889 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1890 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1891 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1892 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1893 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1894 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1895 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1896 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1897 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1898 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1899 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1900 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1901 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1902 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1903 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1904 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1905 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1906 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1907 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1908 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1909 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1910 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1911 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1912 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1913 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1914 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1915 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1916 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1917 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1918 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1919 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1920 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1921 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1922 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1923 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1924 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1925 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1926 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1927 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1928 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1929 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1930 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1931 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1932 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1933 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1934 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1935 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1936 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1937 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1938 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1939 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1940 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1941 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1942 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1943 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1944 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1945 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1946 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1947 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1948 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1949 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1950 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1951 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1952 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1953 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1954 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1955 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1956 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1957 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1958 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1959 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1960 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1961 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1962 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1963 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1964 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1965 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1966 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1967 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1968 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1969 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1970 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1971 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1972 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1973 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1974 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1975 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1976 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1977 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1978 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1979 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1980 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1981 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1982 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1983 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1984 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1985 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1986 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1987 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1988 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1989 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1990 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1991 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1992 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1993 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1994 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1995 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1996 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1997 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1998 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X1999 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2000 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2001 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2002 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2003 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2004 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2005 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2006 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2007 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2008 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2009 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2010 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2011 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2012 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2013 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2014 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2015 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2016 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2017 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2018 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2019 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2020 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2021 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2022 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2023 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2024 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2025 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2026 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2027 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2028 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2029 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2030 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2031 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2032 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2033 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2034 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2035 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2036 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2037 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2038 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2039 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2040 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2041 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2042 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2043 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2044 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2045 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2046 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		X2047 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		
		samples_ready : IN STD_LOGIC := '0';	-- sampler has 2048 samples ready, connected to fft_peripheral pin
		fft_finished : OUT STD_LOGIC := '0';	-- the system is idle / can receive data
		-- clk_in : IN STD_LOGIC;
		
		-- sig_next : OUT STD_LOGIC := '0';
		shift_out0 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000" ;
		shift_out1 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000" ;
		shift_out2 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000" ;
		shift_out3 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000" ;
		shift_out4 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000" ;
		shift_out5 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000" ;
		shift_out6 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000" ;
		shift_out7 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000" ;
		shift_out8 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000" ;
		shift_out9 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000" ;
		shift_out10 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000" ;
		shift_out11 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000" ;
		shift_out12 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000" ;
		shift_out13 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000" ;
		shift_out14 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000" ;
		shift_out15 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000" );
	END COMPONENT;	--c_2048to16x128_shifter
	
	COMPONENT convert2spectrum
		PORT(
		-- R is real and I is imaginary
		X0R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := (others => '0');
		X0I: IN STD_LOGIC_VECTOR(9 DOWNTO 0) := (others => '0');
		X1R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := (others => '0');
		X1I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := (others => '0');
		X2R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := (others => '0');
		X2I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X3R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X3I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X4R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X4I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X5R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X5I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X6R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X6I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X7R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X7I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X8R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X8I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X9R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X9I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X10R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X10I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X11R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X11I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X12R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X12I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X13R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X13I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X14R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X14I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X15R : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X15I : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
	
		V0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
		V1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
		V2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
		V3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
		V4 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
		V5 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
		V6 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
		V7 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
		V8 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
		V9 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
		V10 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
		V11 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
		V12 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
		V13 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
		V14 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
		V15 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
		
		next_bin_set : OUT STD_LOGIC := '0'; -- signal receiving end new bin set data available.
		incoming128set : IN STD_LOGIC := '0'; -- 128 sets of 16 sample incoming
		clk_in : IN STD_LOGIC := '0';
		
		converting : OUT STD_LOGIC := '0');
	END COMPONENT; -- c_10bit2char_vga_H256
	
	BEGIN
		dft_top0 : dft_top
		PORT MAP(
		);
		
		c_2048to16x128_shifter0 : c_2048to16x128_shifter
		PORT MAP(
			X0 <= X0;
		X1 <= X1;
		X2 <= X2;
		X3 <= X3;
		X4 <= X4;
		X5 <= X5;
		X6 <= X6;
		X7 <= X7;
		X8 <= X8;
		X9 <= X9;
		X10 <= X10;
		X11 <= X11;
		X12 <= X12;
		X13 <= X13;
		X14 <= X14;
		X15 <= X15;
		X16 <= X16;
		X17 <= X17;
		X18 <= X18;
		X19 <= X19;
		X20 <= X20;
		X21 <= X21;
		X22 <= X22;
		X23 <= X23;
		X24 <= X24;
		X25 <= X25;
		X26 <= X26;
		X27 <= X27;
		X28 <= X28;
		X29 <= X29;
		X30 <= X30;
		X31 <= X31;
		X32 <= X32;
		X33 <= X33;
		X34 <= X34;
		X35 <= X35;
		X36 <= X36;
		X37 <= X37;
		X38 <= X38;
		X39 <= X39;
		X40 <= X40;
		X41 <= X41;
		X42 <= X42;
		X43 <= X43;
		X44 <= X44;
		X45 <= X45;
		X46 <= X46;
		X47 <= X47;
		X48 <= X48;
		X49 <= X49;
		X50 <= X50;
		X51 <= X51;
		X52 <= X52;
		X53 <= X53;
		X54 <= X54;
		X55 <= X55;
		X56 <= X56;
		X57 <= X57;
		X58 <= X58;
		X59 <= X59;
		X60 <= X60;
		X61 <= X61;
		X62 <= X62;
		X63 <= X63;
		X64 <= X64;
		X65 <= X65;
		X66 <= X66;
		X67 <= X67;
		X68 <= X68;
		X69 <= X69;
		X70 <= X70;
		X71 <= X71;
		X72 <= X72;
		X73 <= X73;
		X74 <= X74;
		X75 <= X75;
		X76 <= X76;
		X77 <= X77;
		X78 <= X78;
		X79 <= X79;
		X80 <= X80;
		X81 <= X81;
		X82 <= X82;
		X83 <= X83;
		X84 <= X84;
		X85 <= X85;
		X86 <= X86;
		X87 <= X87;
		X88 <= X88;
		X89 <= X89;
		X90 <= X90;
		X91 <= X91;
		X92 <= X92;
		X93 <= X93;
		X94 <= X94;
		X95 <= X95;
		X96 <= X96;
		X97 <= X97;
		X98 <= X98;
		X99 <= X99;
		X100 <= X100;
		X101 <= X101;
		X102 <= X102;
		X103 <= X103;
		X104 <= X104;
		X105 <= X105;
		X106 <= X106;
		X107 <= X107;
		X108 <= X108;
		X109 <= X109;
		X110 <= X110;
		X111 <= X111;
		X112 <= X112;
		X113 <= X113;
		X114 <= X114;
		X115 <= X115;
		X116 <= X116;
		X117 <= X117;
		X118 <= X118;
		X119 <= X119;
		X120 <= X120;
		X121 <= X121;
		X122 <= X122;
		X123 <= X123;
		X124 <= X124;
		X125 <= X125;
		X126 <= X126;
		X127 <= X127;
		X128 <= X128;
		X129 <= X129;
		X130 <= X130;
		X131 <= X131;
		X132 <= X132;
		X133 <= X133;
		X134 <= X134;
		X135 <= X135;
		X136 <= X136;
		X137 <= X137;
		X138 <= X138;
		X139 <= X139;
		X140 <= X140;
		X141 <= X141;
		X142 <= X142;
		X143 <= X143;
		X144 <= X144;
		X145 <= X145;
		X146 <= X146;
		X147 <= X147;
		X148 <= X148;
		X149 <= X149;
		X150 <= X150;
		X151 <= X151;
		X152 <= X152;
		X153 <= X153;
		X154 <= X154;
		X155 <= X155;
		X156 <= X156;
		X157 <= X157;
		X158 <= X158;
		X159 <= X159;
		X160 <= X160;
		X161 <= X161;
		X162 <= X162;
		X163 <= X163;
		X164 <= X164;
		X165 <= X165;
		X166 <= X166;
		X167 <= X167;
		X168 <= X168;
		X169 <= X169;
		X170 <= X170;
		X171 <= X171;
		X172 <= X172;
		X173 <= X173;
		X174 <= X174;
		X175 <= X175;
		X176 <= X176;
		X177 <= X177;
		X178 <= X178;
		X179 <= X179;
		X180 <= X180;
		X181 <= X181;
		X182 <= X182;
		X183 <= X183;
		X184 <= X184;
		X185 <= X185;
		X186 <= X186;
		X187 <= X187;
		X188 <= X188;
		X189 <= X189;
		X190 <= X190;
		X191 <= X191;
		X192 <= X192;
		X193 <= X193;
		X194 <= X194;
		X195 <= X195;
		X196 <= X196;
		X197 <= X197;
		X198 <= X198;
		X199 <= X199;
		X200 <= X200;
		X201 <= X201;
		X202 <= X202;
		X203 <= X203;
		X204 <= X204;
		X205 <= X205;
		X206 <= X206;
		X207 <= X207;
		X208 <= X208;
		X209 <= X209;
		X210 <= X210;
		X211 <= X211;
		X212 <= X212;
		X213 <= X213;
		X214 <= X214;
		X215 <= X215;
		X216 <= X216;
		X217 <= X217;
		X218 <= X218;
		X219 <= X219;
		X220 <= X220;
		X221 <= X221;
		X222 <= X222;
		X223 <= X223;
		X224 <= X224;
		X225 <= X225;
		X226 <= X226;
		X227 <= X227;
		X228 <= X228;
		X229 <= X229;
		X230 <= X230;
		X231 <= X231;
		X232 <= X232;
		X233 <= X233;
		X234 <= X234;
		X235 <= X235;
		X236 <= X236;
		X237 <= X237;
		X238 <= X238;
		X239 <= X239;
		X240 <= X240;
		X241 <= X241;
		X242 <= X242;
		X243 <= X243;
		X244 <= X244;
		X245 <= X245;
		X246 <= X246;
		X247 <= X247;
		X248 <= X248;
		X249 <= X249;
		X250 <= X250;
		X251 <= X251;
		X252 <= X252;
		X253 <= X253;
		X254 <= X254;
		X255 <= X255;
		X256 <= X256;
		X257 <= X257;
		X258 <= X258;
		X259 <= X259;
		X260 <= X260;
		X261 <= X261;
		X262 <= X262;
		X263 <= X263;
		X264 <= X264;
		X265 <= X265;
		X266 <= X266;
		X267 <= X267;
		X268 <= X268;
		X269 <= X269;
		X270 <= X270;
		X271 <= X271;
		X272 <= X272;
		X273 <= X273;
		X274 <= X274;
		X275 <= X275;
		X276 <= X276;
		X277 <= X277;
		X278 <= X278;
		X279 <= X279;
		X280 <= X280;
		X281 <= X281;
		X282 <= X282;
		X283 <= X283;
		X284 <= X284;
		X285 <= X285;
		X286 <= X286;
		X287 <= X287;
		X288 <= X288;
		X289 <= X289;
		X290 <= X290;
		X291 <= X291;
		X292 <= X292;
		X293 <= X293;
		X294 <= X294;
		X295 <= X295;
		X296 <= X296;
		X297 <= X297;
		X298 <= X298;
		X299 <= X299;
		X300 <= X300;
		X301 <= X301;
		X302 <= X302;
		X303 <= X303;
		X304 <= X304;
		X305 <= X305;
		X306 <= X306;
		X307 <= X307;
		X308 <= X308;
		X309 <= X309;
		X310 <= X310;
		X311 <= X311;
		X312 <= X312;
		X313 <= X313;
		X314 <= X314;
		X315 <= X315;
		X316 <= X316;
		X317 <= X317;
		X318 <= X318;
		X319 <= X319;
		X320 <= X320;
		X321 <= X321;
		X322 <= X322;
		X323 <= X323;
		X324 <= X324;
		X325 <= X325;
		X326 <= X326;
		X327 <= X327;
		X328 <= X328;
		X329 <= X329;
		X330 <= X330;
		X331 <= X331;
		X332 <= X332;
		X333 <= X333;
		X334 <= X334;
		X335 <= X335;
		X336 <= X336;
		X337 <= X337;
		X338 <= X338;
		X339 <= X339;
		X340 <= X340;
		X341 <= X341;
		X342 <= X342;
		X343 <= X343;
		X344 <= X344;
		X345 <= X345;
		X346 <= X346;
		X347 <= X347;
		X348 <= X348;
		X349 <= X349;
		X350 <= X350;
		X351 <= X351;
		X352 <= X352;
		X353 <= X353;
		X354 <= X354;
		X355 <= X355;
		X356 <= X356;
		X357 <= X357;
		X358 <= X358;
		X359 <= X359;
		X360 <= X360;
		X361 <= X361;
		X362 <= X362;
		X363 <= X363;
		X364 <= X364;
		X365 <= X365;
		X366 <= X366;
		X367 <= X367;
		X368 <= X368;
		X369 <= X369;
		X370 <= X370;
		X371 <= X371;
		X372 <= X372;
		X373 <= X373;
		X374 <= X374;
		X375 <= X375;
		X376 <= X376;
		X377 <= X377;
		X378 <= X378;
		X379 <= X379;
		X380 <= X380;
		X381 <= X381;
		X382 <= X382;
		X383 <= X383;
		X384 <= X384;
		X385 <= X385;
		X386 <= X386;
		X387 <= X387;
		X388 <= X388;
		X389 <= X389;
		X390 <= X390;
		X391 <= X391;
		X392 <= X392;
		X393 <= X393;
		X394 <= X394;
		X395 <= X395;
		X396 <= X396;
		X397 <= X397;
		X398 <= X398;
		X399 <= X399;
		X400 <= X400;
		X401 <= X401;
		X402 <= X402;
		X403 <= X403;
		X404 <= X404;
		X405 <= X405;
		X406 <= X406;
		X407 <= X407;
		X408 <= X408;
		X409 <= X409;
		X410 <= X410;
		X411 <= X411;
		X412 <= X412;
		X413 <= X413;
		X414 <= X414;
		X415 <= X415;
		X416 <= X416;
		X417 <= X417;
		X418 <= X418;
		X419 <= X419;
		X420 <= X420;
		X421 <= X421;
		X422 <= X422;
		X423 <= X423;
		X424 <= X424;
		X425 <= X425;
		X426 <= X426;
		X427 <= X427;
		X428 <= X428;
		X429 <= X429;
		X430 <= X430;
		X431 <= X431;
		X432 <= X432;
		X433 <= X433;
		X434 <= X434;
		X435 <= X435;
		X436 <= X436;
		X437 <= X437;
		X438 <= X438;
		X439 <= X439;
		X440 <= X440;
		X441 <= X441;
		X442 <= X442;
		X443 <= X443;
		X444 <= X444;
		X445 <= X445;
		X446 <= X446;
		X447 <= X447;
		X448 <= X448;
		X449 <= X449;
		X450 <= X450;
		X451 <= X451;
		X452 <= X452;
		X453 <= X453;
		X454 <= X454;
		X455 <= X455;
		X456 <= X456;
		X457 <= X457;
		X458 <= X458;
		X459 <= X459;
		X460 <= X460;
		X461 <= X461;
		X462 <= X462;
		X463 <= X463;
		X464 <= X464;
		X465 <= X465;
		X466 <= X466;
		X467 <= X467;
		X468 <= X468;
		X469 <= X469;
		X470 <= X470;
		X471 <= X471;
		X472 <= X472;
		X473 <= X473;
		X474 <= X474;
		X475 <= X475;
		X476 <= X476;
		X477 <= X477;
		X478 <= X478;
		X479 <= X479;
		X480 <= X480;
		X481 <= X481;
		X482 <= X482;
		X483 <= X483;
		X484 <= X484;
		X485 <= X485;
		X486 <= X486;
		X487 <= X487;
		X488 <= X488;
		X489 <= X489;
		X490 <= X490;
		X491 <= X491;
		X492 <= X492;
		X493 <= X493;
		X494 <= X494;
		X495 <= X495;
		X496 <= X496;
		X497 <= X497;
		X498 <= X498;
		X499 <= X499;
		X500 <= X500;
		X501 <= X501;
		X502 <= X502;
		X503 <= X503;
		X504 <= X504;
		X505 <= X505;
		X506 <= X506;
		X507 <= X507;
		X508 <= X508;
		X509 <= X509;
		X510 <= X510;
		X511 <= X511;
		X512 <= X512;
		X513 <= X513;
		X514 <= X514;
		X515 <= X515;
		X516 <= X516;
		X517 <= X517;
		X518 <= X518;
		X519 <= X519;
		X520 <= X520;
		X521 <= X521;
		X522 <= X522;
		X523 <= X523;
		X524 <= X524;
		X525 <= X525;
		X526 <= X526;
		X527 <= X527;
		X528 <= X528;
		X529 <= X529;
		X530 <= X530;
		X531 <= X531;
		X532 <= X532;
		X533 <= X533;
		X534 <= X534;
		X535 <= X535;
		X536 <= X536;
		X537 <= X537;
		X538 <= X538;
		X539 <= X539;
		X540 <= X540;
		X541 <= X541;
		X542 <= X542;
		X543 <= X543;
		X544 <= X544;
		X545 <= X545;
		X546 <= X546;
		X547 <= X547;
		X548 <= X548;
		X549 <= X549;
		X550 <= X550;
		X551 <= X551;
		X552 <= X552;
		X553 <= X553;
		X554 <= X554;
		X555 <= X555;
		X556 <= X556;
		X557 <= X557;
		X558 <= X558;
		X559 <= X559;
		X560 <= X560;
		X561 <= X561;
		X562 <= X562;
		X563 <= X563;
		X564 <= X564;
		X565 <= X565;
		X566 <= X566;
		X567 <= X567;
		X568 <= X568;
		X569 <= X569;
		X570 <= X570;
		X571 <= X571;
		X572 <= X572;
		X573 <= X573;
		X574 <= X574;
		X575 <= X575;
		X576 <= X576;
		X577 <= X577;
		X578 <= X578;
		X579 <= X579;
		X580 <= X580;
		X581 <= X581;
		X582 <= X582;
		X583 <= X583;
		X584 <= X584;
		X585 <= X585;
		X586 <= X586;
		X587 <= X587;
		X588 <= X588;
		X589 <= X589;
		X590 <= X590;
		X591 <= X591;
		X592 <= X592;
		X593 <= X593;
		X594 <= X594;
		X595 <= X595;
		X596 <= X596;
		X597 <= X597;
		X598 <= X598;
		X599 <= X599;
		X600 <= X600;
		X601 <= X601;
		X602 <= X602;
		X603 <= X603;
		X604 <= X604;
		X605 <= X605;
		X606 <= X606;
		X607 <= X607;
		X608 <= X608;
		X609 <= X609;
		X610 <= X610;
		X611 <= X611;
		X612 <= X612;
		X613 <= X613;
		X614 <= X614;
		X615 <= X615;
		X616 <= X616;
		X617 <= X617;
		X618 <= X618;
		X619 <= X619;
		X620 <= X620;
		X621 <= X621;
		X622 <= X622;
		X623 <= X623;
		X624 <= X624;
		X625 <= X625;
		X626 <= X626;
		X627 <= X627;
		X628 <= X628;
		X629 <= X629;
		X630 <= X630;
		X631 <= X631;
		X632 <= X632;
		X633 <= X633;
		X634 <= X634;
		X635 <= X635;
		X636 <= X636;
		X637 <= X637;
		X638 <= X638;
		X639 <= X639;
		X640 <= X640;
		X641 <= X641;
		X642 <= X642;
		X643 <= X643;
		X644 <= X644;
		X645 <= X645;
		X646 <= X646;
		X647 <= X647;
		X648 <= X648;
		X649 <= X649;
		X650 <= X650;
		X651 <= X651;
		X652 <= X652;
		X653 <= X653;
		X654 <= X654;
		X655 <= X655;
		X656 <= X656;
		X657 <= X657;
		X658 <= X658;
		X659 <= X659;
		X660 <= X660;
		X661 <= X661;
		X662 <= X662;
		X663 <= X663;
		X664 <= X664;
		X665 <= X665;
		X666 <= X666;
		X667 <= X667;
		X668 <= X668;
		X669 <= X669;
		X670 <= X670;
		X671 <= X671;
		X672 <= X672;
		X673 <= X673;
		X674 <= X674;
		X675 <= X675;
		X676 <= X676;
		X677 <= X677;
		X678 <= X678;
		X679 <= X679;
		X680 <= X680;
		X681 <= X681;
		X682 <= X682;
		X683 <= X683;
		X684 <= X684;
		X685 <= X685;
		X686 <= X686;
		X687 <= X687;
		X688 <= X688;
		X689 <= X689;
		X690 <= X690;
		X691 <= X691;
		X692 <= X692;
		X693 <= X693;
		X694 <= X694;
		X695 <= X695;
		X696 <= X696;
		X697 <= X697;
		X698 <= X698;
		X699 <= X699;
		X700 <= X700;
		X701 <= X701;
		X702 <= X702;
		X703 <= X703;
		X704 <= X704;
		X705 <= X705;
		X706 <= X706;
		X707 <= X707;
		X708 <= X708;
		X709 <= X709;
		X710 <= X710;
		X711 <= X711;
		X712 <= X712;
		X713 <= X713;
		X714 <= X714;
		X715 <= X715;
		X716 <= X716;
		X717 <= X717;
		X718 <= X718;
		X719 <= X719;
		X720 <= X720;
		X721 <= X721;
		X722 <= X722;
		X723 <= X723;
		X724 <= X724;
		X725 <= X725;
		X726 <= X726;
		X727 <= X727;
		X728 <= X728;
		X729 <= X729;
		X730 <= X730;
		X731 <= X731;
		X732 <= X732;
		X733 <= X733;
		X734 <= X734;
		X735 <= X735;
		X736 <= X736;
		X737 <= X737;
		X738 <= X738;
		X739 <= X739;
		X740 <= X740;
		X741 <= X741;
		X742 <= X742;
		X743 <= X743;
		X744 <= X744;
		X745 <= X745;
		X746 <= X746;
		X747 <= X747;
		X748 <= X748;
		X749 <= X749;
		X750 <= X750;
		X751 <= X751;
		X752 <= X752;
		X753 <= X753;
		X754 <= X754;
		X755 <= X755;
		X756 <= X756;
		X757 <= X757;
		X758 <= X758;
		X759 <= X759;
		X760 <= X760;
		X761 <= X761;
		X762 <= X762;
		X763 <= X763;
		X764 <= X764;
		X765 <= X765;
		X766 <= X766;
		X767 <= X767;
		X768 <= X768;
		X769 <= X769;
		X770 <= X770;
		X771 <= X771;
		X772 <= X772;
		X773 <= X773;
		X774 <= X774;
		X775 <= X775;
		X776 <= X776;
		X777 <= X777;
		X778 <= X778;
		X779 <= X779;
		X780 <= X780;
		X781 <= X781;
		X782 <= X782;
		X783 <= X783;
		X784 <= X784;
		X785 <= X785;
		X786 <= X786;
		X787 <= X787;
		X788 <= X788;
		X789 <= X789;
		X790 <= X790;
		X791 <= X791;
		X792 <= X792;
		X793 <= X793;
		X794 <= X794;
		X795 <= X795;
		X796 <= X796;
		X797 <= X797;
		X798 <= X798;
		X799 <= X799;
		X800 <= X800;
		X801 <= X801;
		X802 <= X802;
		X803 <= X803;
		X804 <= X804;
		X805 <= X805;
		X806 <= X806;
		X807 <= X807;
		X808 <= X808;
		X809 <= X809;
		X810 <= X810;
		X811 <= X811;
		X812 <= X812;
		X813 <= X813;
		X814 <= X814;
		X815 <= X815;
		X816 <= X816;
		X817 <= X817;
		X818 <= X818;
		X819 <= X819;
		X820 <= X820;
		X821 <= X821;
		X822 <= X822;
		X823 <= X823;
		X824 <= X824;
		X825 <= X825;
		X826 <= X826;
		X827 <= X827;
		X828 <= X828;
		X829 <= X829;
		X830 <= X830;
		X831 <= X831;
		X832 <= X832;
		X833 <= X833;
		X834 <= X834;
		X835 <= X835;
		X836 <= X836;
		X837 <= X837;
		X838 <= X838;
		X839 <= X839;
		X840 <= X840;
		X841 <= X841;
		X842 <= X842;
		X843 <= X843;
		X844 <= X844;
		X845 <= X845;
		X846 <= X846;
		X847 <= X847;
		X848 <= X848;
		X849 <= X849;
		X850 <= X850;
		X851 <= X851;
		X852 <= X852;
		X853 <= X853;
		X854 <= X854;
		X855 <= X855;
		X856 <= X856;
		X857 <= X857;
		X858 <= X858;
		X859 <= X859;
		X860 <= X860;
		X861 <= X861;
		X862 <= X862;
		X863 <= X863;
		X864 <= X864;
		X865 <= X865;
		X866 <= X866;
		X867 <= X867;
		X868 <= X868;
		X869 <= X869;
		X870 <= X870;
		X871 <= X871;
		X872 <= X872;
		X873 <= X873;
		X874 <= X874;
		X875 <= X875;
		X876 <= X876;
		X877 <= X877;
		X878 <= X878;
		X879 <= X879;
		X880 <= X880;
		X881 <= X881;
		X882 <= X882;
		X883 <= X883;
		X884 <= X884;
		X885 <= X885;
		X886 <= X886;
		X887 <= X887;
		X888 <= X888;
		X889 <= X889;
		X890 <= X890;
		X891 <= X891;
		X892 <= X892;
		X893 <= X893;
		X894 <= X894;
		X895 <= X895;
		X896 <= X896;
		X897 <= X897;
		X898 <= X898;
		X899 <= X899;
		X900 <= X900;
		X901 <= X901;
		X902 <= X902;
		X903 <= X903;
		X904 <= X904;
		X905 <= X905;
		X906 <= X906;
		X907 <= X907;
		X908 <= X908;
		X909 <= X909;
		X910 <= X910;
		X911 <= X911;
		X912 <= X912;
		X913 <= X913;
		X914 <= X914;
		X915 <= X915;
		X916 <= X916;
		X917 <= X917;
		X918 <= X918;
		X919 <= X919;
		X920 <= X920;
		X921 <= X921;
		X922 <= X922;
		X923 <= X923;
		X924 <= X924;
		X925 <= X925;
		X926 <= X926;
		X927 <= X927;
		X928 <= X928;
		X929 <= X929;
		X930 <= X930;
		X931 <= X931;
		X932 <= X932;
		X933 <= X933;
		X934 <= X934;
		X935 <= X935;
		X936 <= X936;
		X937 <= X937;
		X938 <= X938;
		X939 <= X939;
		X940 <= X940;
		X941 <= X941;
		X942 <= X942;
		X943 <= X943;
		X944 <= X944;
		X945 <= X945;
		X946 <= X946;
		X947 <= X947;
		X948 <= X948;
		X949 <= X949;
		X950 <= X950;
		X951 <= X951;
		X952 <= X952;
		X953 <= X953;
		X954 <= X954;
		X955 <= X955;
		X956 <= X956;
		X957 <= X957;
		X958 <= X958;
		X959 <= X959;
		X960 <= X960;
		X961 <= X961;
		X962 <= X962;
		X963 <= X963;
		X964 <= X964;
		X965 <= X965;
		X966 <= X966;
		X967 <= X967;
		X968 <= X968;
		X969 <= X969;
		X970 <= X970;
		X971 <= X971;
		X972 <= X972;
		X973 <= X973;
		X974 <= X974;
		X975 <= X975;
		X976 <= X976;
		X977 <= X977;
		X978 <= X978;
		X979 <= X979;
		X980 <= X980;
		X981 <= X981;
		X982 <= X982;
		X983 <= X983;
		X984 <= X984;
		X985 <= X985;
		X986 <= X986;
		X987 <= X987;
		X988 <= X988;
		X989 <= X989;
		X990 <= X990;
		X991 <= X991;
		X992 <= X992;
		X993 <= X993;
		X994 <= X994;
		X995 <= X995;
		X996 <= X996;
		X997 <= X997;
		X998 <= X998;
		X999 <= X999;
		X1000 <= X1000;
		X1001 <= X1001;
		X1002 <= X1002;
		X1003 <= X1003;
		X1004 <= X1004;
		X1005 <= X1005;
		X1006 <= X1006;
		X1007 <= X1007;
		X1008 <= X1008;
		X1009 <= X1009;
		X1010 <= X1010;
		X1011 <= X1011;
		X1012 <= X1012;
		X1013 <= X1013;
		X1014 <= X1014;
		X1015 <= X1015;
		X1016 <= X1016;
		X1017 <= X1017;
		X1018 <= X1018;
		X1019 <= X1019;
		X1020 <= X1020;
		X1021 <= X1021;
		X1022 <= X1022;
		X1023 <= X1023;
		X1024 <= X1024;
		X1025 <= X1025;
		X1026 <= X1026;
		X1027 <= X1027;
		X1028 <= X1028;
		X1029 <= X1029;
		X1030 <= X1030;
		X1031 <= X1031;
		X1032 <= X1032;
		X1033 <= X1033;
		X1034 <= X1034;
		X1035 <= X1035;
		X1036 <= X1036;
		X1037 <= X1037;
		X1038 <= X1038;
		X1039 <= X1039;
		X1040 <= X1040;
		X1041 <= X1041;
		X1042 <= X1042;
		X1043 <= X1043;
		X1044 <= X1044;
		X1045 <= X1045;
		X1046 <= X1046;
		X1047 <= X1047;
		X1048 <= X1048;
		X1049 <= X1049;
		X1050 <= X1050;
		X1051 <= X1051;
		X1052 <= X1052;
		X1053 <= X1053;
		X1054 <= X1054;
		X1055 <= X1055;
		X1056 <= X1056;
		X1057 <= X1057;
		X1058 <= X1058;
		X1059 <= X1059;
		X1060 <= X1060;
		X1061 <= X1061;
		X1062 <= X1062;
		X1063 <= X1063;
		X1064 <= X1064;
		X1065 <= X1065;
		X1066 <= X1066;
		X1067 <= X1067;
		X1068 <= X1068;
		X1069 <= X1069;
		X1070 <= X1070;
		X1071 <= X1071;
		X1072 <= X1072;
		X1073 <= X1073;
		X1074 <= X1074;
		X1075 <= X1075;
		X1076 <= X1076;
		X1077 <= X1077;
		X1078 <= X1078;
		X1079 <= X1079;
		X1080 <= X1080;
		X1081 <= X1081;
		X1082 <= X1082;
		X1083 <= X1083;
		X1084 <= X1084;
		X1085 <= X1085;
		X1086 <= X1086;
		X1087 <= X1087;
		X1088 <= X1088;
		X1089 <= X1089;
		X1090 <= X1090;
		X1091 <= X1091;
		X1092 <= X1092;
		X1093 <= X1093;
		X1094 <= X1094;
		X1095 <= X1095;
		X1096 <= X1096;
		X1097 <= X1097;
		X1098 <= X1098;
		X1099 <= X1099;
		X1100 <= X1100;
		X1101 <= X1101;
		X1102 <= X1102;
		X1103 <= X1103;
		X1104 <= X1104;
		X1105 <= X1105;
		X1106 <= X1106;
		X1107 <= X1107;
		X1108 <= X1108;
		X1109 <= X1109;
		X1110 <= X1110;
		X1111 <= X1111;
		X1112 <= X1112;
		X1113 <= X1113;
		X1114 <= X1114;
		X1115 <= X1115;
		X1116 <= X1116;
		X1117 <= X1117;
		X1118 <= X1118;
		X1119 <= X1119;
		X1120 <= X1120;
		X1121 <= X1121;
		X1122 <= X1122;
		X1123 <= X1123;
		X1124 <= X1124;
		X1125 <= X1125;
		X1126 <= X1126;
		X1127 <= X1127;
		X1128 <= X1128;
		X1129 <= X1129;
		X1130 <= X1130;
		X1131 <= X1131;
		X1132 <= X1132;
		X1133 <= X1133;
		X1134 <= X1134;
		X1135 <= X1135;
		X1136 <= X1136;
		X1137 <= X1137;
		X1138 <= X1138;
		X1139 <= X1139;
		X1140 <= X1140;
		X1141 <= X1141;
		X1142 <= X1142;
		X1143 <= X1143;
		X1144 <= X1144;
		X1145 <= X1145;
		X1146 <= X1146;
		X1147 <= X1147;
		X1148 <= X1148;
		X1149 <= X1149;
		X1150 <= X1150;
		X1151 <= X1151;
		X1152 <= X1152;
		X1153 <= X1153;
		X1154 <= X1154;
		X1155 <= X1155;
		X1156 <= X1156;
		X1157 <= X1157;
		X1158 <= X1158;
		X1159 <= X1159;
		X1160 <= X1160;
		X1161 <= X1161;
		X1162 <= X1162;
		X1163 <= X1163;
		X1164 <= X1164;
		X1165 <= X1165;
		X1166 <= X1166;
		X1167 <= X1167;
		X1168 <= X1168;
		X1169 <= X1169;
		X1170 <= X1170;
		X1171 <= X1171;
		X1172 <= X1172;
		X1173 <= X1173;
		X1174 <= X1174;
		X1175 <= X1175;
		X1176 <= X1176;
		X1177 <= X1177;
		X1178 <= X1178;
		X1179 <= X1179;
		X1180 <= X1180;
		X1181 <= X1181;
		X1182 <= X1182;
		X1183 <= X1183;
		X1184 <= X1184;
		X1185 <= X1185;
		X1186 <= X1186;
		X1187 <= X1187;
		X1188 <= X1188;
		X1189 <= X1189;
		X1190 <= X1190;
		X1191 <= X1191;
		X1192 <= X1192;
		X1193 <= X1193;
		X1194 <= X1194;
		X1195 <= X1195;
		X1196 <= X1196;
		X1197 <= X1197;
		X1198 <= X1198;
		X1199 <= X1199;
		X1200 <= X1200;
		X1201 <= X1201;
		X1202 <= X1202;
		X1203 <= X1203;
		X1204 <= X1204;
		X1205 <= X1205;
		X1206 <= X1206;
		X1207 <= X1207;
		X1208 <= X1208;
		X1209 <= X1209;
		X1210 <= X1210;
		X1211 <= X1211;
		X1212 <= X1212;
		X1213 <= X1213;
		X1214 <= X1214;
		X1215 <= X1215;
		X1216 <= X1216;
		X1217 <= X1217;
		X1218 <= X1218;
		X1219 <= X1219;
		X1220 <= X1220;
		X1221 <= X1221;
		X1222 <= X1222;
		X1223 <= X1223;
		X1224 <= X1224;
		X1225 <= X1225;
		X1226 <= X1226;
		X1227 <= X1227;
		X1228 <= X1228;
		X1229 <= X1229;
		X1230 <= X1230;
		X1231 <= X1231;
		X1232 <= X1232;
		X1233 <= X1233;
		X1234 <= X1234;
		X1235 <= X1235;
		X1236 <= X1236;
		X1237 <= X1237;
		X1238 <= X1238;
		X1239 <= X1239;
		X1240 <= X1240;
		X1241 <= X1241;
		X1242 <= X1242;
		X1243 <= X1243;
		X1244 <= X1244;
		X1245 <= X1245;
		X1246 <= X1246;
		X1247 <= X1247;
		X1248 <= X1248;
		X1249 <= X1249;
		X1250 <= X1250;
		X1251 <= X1251;
		X1252 <= X1252;
		X1253 <= X1253;
		X1254 <= X1254;
		X1255 <= X1255;
		X1256 <= X1256;
		X1257 <= X1257;
		X1258 <= X1258;
		X1259 <= X1259;
		X1260 <= X1260;
		X1261 <= X1261;
		X1262 <= X1262;
		X1263 <= X1263;
		X1264 <= X1264;
		X1265 <= X1265;
		X1266 <= X1266;
		X1267 <= X1267;
		X1268 <= X1268;
		X1269 <= X1269;
		X1270 <= X1270;
		X1271 <= X1271;
		X1272 <= X1272;
		X1273 <= X1273;
		X1274 <= X1274;
		X1275 <= X1275;
		X1276 <= X1276;
		X1277 <= X1277;
		X1278 <= X1278;
		X1279 <= X1279;
		X1280 <= X1280;
		X1281 <= X1281;
		X1282 <= X1282;
		X1283 <= X1283;
		X1284 <= X1284;
		X1285 <= X1285;
		X1286 <= X1286;
		X1287 <= X1287;
		X1288 <= X1288;
		X1289 <= X1289;
		X1290 <= X1290;
		X1291 <= X1291;
		X1292 <= X1292;
		X1293 <= X1293;
		X1294 <= X1294;
		X1295 <= X1295;
		X1296 <= X1296;
		X1297 <= X1297;
		X1298 <= X1298;
		X1299 <= X1299;
		X1300 <= X1300;
		X1301 <= X1301;
		X1302 <= X1302;
		X1303 <= X1303;
		X1304 <= X1304;
		X1305 <= X1305;
		X1306 <= X1306;
		X1307 <= X1307;
		X1308 <= X1308;
		X1309 <= X1309;
		X1310 <= X1310;
		X1311 <= X1311;
		X1312 <= X1312;
		X1313 <= X1313;
		X1314 <= X1314;
		X1315 <= X1315;
		X1316 <= X1316;
		X1317 <= X1317;
		X1318 <= X1318;
		X1319 <= X1319;
		X1320 <= X1320;
		X1321 <= X1321;
		X1322 <= X1322;
		X1323 <= X1323;
		X1324 <= X1324;
		X1325 <= X1325;
		X1326 <= X1326;
		X1327 <= X1327;
		X1328 <= X1328;
		X1329 <= X1329;
		X1330 <= X1330;
		X1331 <= X1331;
		X1332 <= X1332;
		X1333 <= X1333;
		X1334 <= X1334;
		X1335 <= X1335;
		X1336 <= X1336;
		X1337 <= X1337;
		X1338 <= X1338;
		X1339 <= X1339;
		X1340 <= X1340;
		X1341 <= X1341;
		X1342 <= X1342;
		X1343 <= X1343;
		X1344 <= X1344;
		X1345 <= X1345;
		X1346 <= X1346;
		X1347 <= X1347;
		X1348 <= X1348;
		X1349 <= X1349;
		X1350 <= X1350;
		X1351 <= X1351;
		X1352 <= X1352;
		X1353 <= X1353;
		X1354 <= X1354;
		X1355 <= X1355;
		X1356 <= X1356;
		X1357 <= X1357;
		X1358 <= X1358;
		X1359 <= X1359;
		X1360 <= X1360;
		X1361 <= X1361;
		X1362 <= X1362;
		X1363 <= X1363;
		X1364 <= X1364;
		X1365 <= X1365;
		X1366 <= X1366;
		X1367 <= X1367;
		X1368 <= X1368;
		X1369 <= X1369;
		X1370 <= X1370;
		X1371 <= X1371;
		X1372 <= X1372;
		X1373 <= X1373;
		X1374 <= X1374;
		X1375 <= X1375;
		X1376 <= X1376;
		X1377 <= X1377;
		X1378 <= X1378;
		X1379 <= X1379;
		X1380 <= X1380;
		X1381 <= X1381;
		X1382 <= X1382;
		X1383 <= X1383;
		X1384 <= X1384;
		X1385 <= X1385;
		X1386 <= X1386;
		X1387 <= X1387;
		X1388 <= X1388;
		X1389 <= X1389;
		X1390 <= X1390;
		X1391 <= X1391;
		X1392 <= X1392;
		X1393 <= X1393;
		X1394 <= X1394;
		X1395 <= X1395;
		X1396 <= X1396;
		X1397 <= X1397;
		X1398 <= X1398;
		X1399 <= X1399;
		X1400 <= X1400;
		X1401 <= X1401;
		X1402 <= X1402;
		X1403 <= X1403;
		X1404 <= X1404;
		X1405 <= X1405;
		X1406 <= X1406;
		X1407 <= X1407;
		X1408 <= X1408;
		X1409 <= X1409;
		X1410 <= X1410;
		X1411 <= X1411;
		X1412 <= X1412;
		X1413 <= X1413;
		X1414 <= X1414;
		X1415 <= X1415;
		X1416 <= X1416;
		X1417 <= X1417;
		X1418 <= X1418;
		X1419 <= X1419;
		X1420 <= X1420;
		X1421 <= X1421;
		X1422 <= X1422;
		X1423 <= X1423;
		X1424 <= X1424;
		X1425 <= X1425;
		X1426 <= X1426;
		X1427 <= X1427;
		X1428 <= X1428;
		X1429 <= X1429;
		X1430 <= X1430;
		X1431 <= X1431;
		X1432 <= X1432;
		X1433 <= X1433;
		X1434 <= X1434;
		X1435 <= X1435;
		X1436 <= X1436;
		X1437 <= X1437;
		X1438 <= X1438;
		X1439 <= X1439;
		X1440 <= X1440;
		X1441 <= X1441;
		X1442 <= X1442;
		X1443 <= X1443;
		X1444 <= X1444;
		X1445 <= X1445;
		X1446 <= X1446;
		X1447 <= X1447;
		X1448 <= X1448;
		X1449 <= X1449;
		X1450 <= X1450;
		X1451 <= X1451;
		X1452 <= X1452;
		X1453 <= X1453;
		X1454 <= X1454;
		X1455 <= X1455;
		X1456 <= X1456;
		X1457 <= X1457;
		X1458 <= X1458;
		X1459 <= X1459;
		X1460 <= X1460;
		X1461 <= X1461;
		X1462 <= X1462;
		X1463 <= X1463;
		X1464 <= X1464;
		X1465 <= X1465;
		X1466 <= X1466;
		X1467 <= X1467;
		X1468 <= X1468;
		X1469 <= X1469;
		X1470 <= X1470;
		X1471 <= X1471;
		X1472 <= X1472;
		X1473 <= X1473;
		X1474 <= X1474;
		X1475 <= X1475;
		X1476 <= X1476;
		X1477 <= X1477;
		X1478 <= X1478;
		X1479 <= X1479;
		X1480 <= X1480;
		X1481 <= X1481;
		X1482 <= X1482;
		X1483 <= X1483;
		X1484 <= X1484;
		X1485 <= X1485;
		X1486 <= X1486;
		X1487 <= X1487;
		X1488 <= X1488;
		X1489 <= X1489;
		X1490 <= X1490;
		X1491 <= X1491;
		X1492 <= X1492;
		X1493 <= X1493;
		X1494 <= X1494;
		X1495 <= X1495;
		X1496 <= X1496;
		X1497 <= X1497;
		X1498 <= X1498;
		X1499 <= X1499;
		X1500 <= X1500;
		X1501 <= X1501;
		X1502 <= X1502;
		X1503 <= X1503;
		X1504 <= X1504;
		X1505 <= X1505;
		X1506 <= X1506;
		X1507 <= X1507;
		X1508 <= X1508;
		X1509 <= X1509;
		X1510 <= X1510;
		X1511 <= X1511;
		X1512 <= X1512;
		X1513 <= X1513;
		X1514 <= X1514;
		X1515 <= X1515;
		X1516 <= X1516;
		X1517 <= X1517;
		X1518 <= X1518;
		X1519 <= X1519;
		X1520 <= X1520;
		X1521 <= X1521;
		X1522 <= X1522;
		X1523 <= X1523;
		X1524 <= X1524;
		X1525 <= X1525;
		X1526 <= X1526;
		X1527 <= X1527;
		X1528 <= X1528;
		X1529 <= X1529;
		X1530 <= X1530;
		X1531 <= X1531;
		X1532 <= X1532;
		X1533 <= X1533;
		X1534 <= X1534;
		X1535 <= X1535;
		X1536 <= X1536;
		X1537 <= X1537;
		X1538 <= X1538;
		X1539 <= X1539;
		X1540 <= X1540;
		X1541 <= X1541;
		X1542 <= X1542;
		X1543 <= X1543;
		X1544 <= X1544;
		X1545 <= X1545;
		X1546 <= X1546;
		X1547 <= X1547;
		X1548 <= X1548;
		X1549 <= X1549;
		X1550 <= X1550;
		X1551 <= X1551;
		X1552 <= X1552;
		X1553 <= X1553;
		X1554 <= X1554;
		X1555 <= X1555;
		X1556 <= X1556;
		X1557 <= X1557;
		X1558 <= X1558;
		X1559 <= X1559;
		X1560 <= X1560;
		X1561 <= X1561;
		X1562 <= X1562;
		X1563 <= X1563;
		X1564 <= X1564;
		X1565 <= X1565;
		X1566 <= X1566;
		X1567 <= X1567;
		X1568 <= X1568;
		X1569 <= X1569;
		X1570 <= X1570;
		X1571 <= X1571;
		X1572 <= X1572;
		X1573 <= X1573;
		X1574 <= X1574;
		X1575 <= X1575;
		X1576 <= X1576;
		X1577 <= X1577;
		X1578 <= X1578;
		X1579 <= X1579;
		X1580 <= X1580;
		X1581 <= X1581;
		X1582 <= X1582;
		X1583 <= X1583;
		X1584 <= X1584;
		X1585 <= X1585;
		X1586 <= X1586;
		X1587 <= X1587;
		X1588 <= X1588;
		X1589 <= X1589;
		X1590 <= X1590;
		X1591 <= X1591;
		X1592 <= X1592;
		X1593 <= X1593;
		X1594 <= X1594;
		X1595 <= X1595;
		X1596 <= X1596;
		X1597 <= X1597;
		X1598 <= X1598;
		X1599 <= X1599;
		X1600 <= X1600;
		X1601 <= X1601;
		X1602 <= X1602;
		X1603 <= X1603;
		X1604 <= X1604;
		X1605 <= X1605;
		X1606 <= X1606;
		X1607 <= X1607;
		X1608 <= X1608;
		X1609 <= X1609;
		X1610 <= X1610;
		X1611 <= X1611;
		X1612 <= X1612;
		X1613 <= X1613;
		X1614 <= X1614;
		X1615 <= X1615;
		X1616 <= X1616;
		X1617 <= X1617;
		X1618 <= X1618;
		X1619 <= X1619;
		X1620 <= X1620;
		X1621 <= X1621;
		X1622 <= X1622;
		X1623 <= X1623;
		X1624 <= X1624;
		X1625 <= X1625;
		X1626 <= X1626;
		X1627 <= X1627;
		X1628 <= X1628;
		X1629 <= X1629;
		X1630 <= X1630;
		X1631 <= X1631;
		X1632 <= X1632;
		X1633 <= X1633;
		X1634 <= X1634;
		X1635 <= X1635;
		X1636 <= X1636;
		X1637 <= X1637;
		X1638 <= X1638;
		X1639 <= X1639;
		X1640 <= X1640;
		X1641 <= X1641;
		X1642 <= X1642;
		X1643 <= X1643;
		X1644 <= X1644;
		X1645 <= X1645;
		X1646 <= X1646;
		X1647 <= X1647;
		X1648 <= X1648;
		X1649 <= X1649;
		X1650 <= X1650;
		X1651 <= X1651;
		X1652 <= X1652;
		X1653 <= X1653;
		X1654 <= X1654;
		X1655 <= X1655;
		X1656 <= X1656;
		X1657 <= X1657;
		X1658 <= X1658;
		X1659 <= X1659;
		X1660 <= X1660;
		X1661 <= X1661;
		X1662 <= X1662;
		X1663 <= X1663;
		X1664 <= X1664;
		X1665 <= X1665;
		X1666 <= X1666;
		X1667 <= X1667;
		X1668 <= X1668;
		X1669 <= X1669;
		X1670 <= X1670;
		X1671 <= X1671;
		X1672 <= X1672;
		X1673 <= X1673;
		X1674 <= X1674;
		X1675 <= X1675;
		X1676 <= X1676;
		X1677 <= X1677;
		X1678 <= X1678;
		X1679 <= X1679;
		X1680 <= X1680;
		X1681 <= X1681;
		X1682 <= X1682;
		X1683 <= X1683;
		X1684 <= X1684;
		X1685 <= X1685;
		X1686 <= X1686;
		X1687 <= X1687;
		X1688 <= X1688;
		X1689 <= X1689;
		X1690 <= X1690;
		X1691 <= X1691;
		X1692 <= X1692;
		X1693 <= X1693;
		X1694 <= X1694;
		X1695 <= X1695;
		X1696 <= X1696;
		X1697 <= X1697;
		X1698 <= X1698;
		X1699 <= X1699;
		X1700 <= X1700;
		X1701 <= X1701;
		X1702 <= X1702;
		X1703 <= X1703;
		X1704 <= X1704;
		X1705 <= X1705;
		X1706 <= X1706;
		X1707 <= X1707;
		X1708 <= X1708;
		X1709 <= X1709;
		X1710 <= X1710;
		X1711 <= X1711;
		X1712 <= X1712;
		X1713 <= X1713;
		X1714 <= X1714;
		X1715 <= X1715;
		X1716 <= X1716;
		X1717 <= X1717;
		X1718 <= X1718;
		X1719 <= X1719;
		X1720 <= X1720;
		X1721 <= X1721;
		X1722 <= X1722;
		X1723 <= X1723;
		X1724 <= X1724;
		X1725 <= X1725;
		X1726 <= X1726;
		X1727 <= X1727;
		X1728 <= X1728;
		X1729 <= X1729;
		X1730 <= X1730;
		X1731 <= X1731;
		X1732 <= X1732;
		X1733 <= X1733;
		X1734 <= X1734;
		X1735 <= X1735;
		X1736 <= X1736;
		X1737 <= X1737;
		X1738 <= X1738;
		X1739 <= X1739;
		X1740 <= X1740;
		X1741 <= X1741;
		X1742 <= X1742;
		X1743 <= X1743;
		X1744 <= X1744;
		X1745 <= X1745;
		X1746 <= X1746;
		X1747 <= X1747;
		X1748 <= X1748;
		X1749 <= X1749;
		X1750 <= X1750;
		X1751 <= X1751;
		X1752 <= X1752;
		X1753 <= X1753;
		X1754 <= X1754;
		X1755 <= X1755;
		X1756 <= X1756;
		X1757 <= X1757;
		X1758 <= X1758;
		X1759 <= X1759;
		X1760 <= X1760;
		X1761 <= X1761;
		X1762 <= X1762;
		X1763 <= X1763;
		X1764 <= X1764;
		X1765 <= X1765;
		X1766 <= X1766;
		X1767 <= X1767;
		X1768 <= X1768;
		X1769 <= X1769;
		X1770 <= X1770;
		X1771 <= X1771;
		X1772 <= X1772;
		X1773 <= X1773;
		X1774 <= X1774;
		X1775 <= X1775;
		X1776 <= X1776;
		X1777 <= X1777;
		X1778 <= X1778;
		X1779 <= X1779;
		X1780 <= X1780;
		X1781 <= X1781;
		X1782 <= X1782;
		X1783 <= X1783;
		X1784 <= X1784;
		X1785 <= X1785;
		X1786 <= X1786;
		X1787 <= X1787;
		X1788 <= X1788;
		X1789 <= X1789;
		X1790 <= X1790;
		X1791 <= X1791;
		X1792 <= X1792;
		X1793 <= X1793;
		X1794 <= X1794;
		X1795 <= X1795;
		X1796 <= X1796;
		X1797 <= X1797;
		X1798 <= X1798;
		X1799 <= X1799;
		X1800 <= X1800;
		X1801 <= X1801;
		X1802 <= X1802;
		X1803 <= X1803;
		X1804 <= X1804;
		X1805 <= X1805;
		X1806 <= X1806;
		X1807 <= X1807;
		X1808 <= X1808;
		X1809 <= X1809;
		X1810 <= X1810;
		X1811 <= X1811;
		X1812 <= X1812;
		X1813 <= X1813;
		X1814 <= X1814;
		X1815 <= X1815;
		X1816 <= X1816;
		X1817 <= X1817;
		X1818 <= X1818;
		X1819 <= X1819;
		X1820 <= X1820;
		X1821 <= X1821;
		X1822 <= X1822;
		X1823 <= X1823;
		X1824 <= X1824;
		X1825 <= X1825;
		X1826 <= X1826;
		X1827 <= X1827;
		X1828 <= X1828;
		X1829 <= X1829;
		X1830 <= X1830;
		X1831 <= X1831;
		X1832 <= X1832;
		X1833 <= X1833;
		X1834 <= X1834;
		X1835 <= X1835;
		X1836 <= X1836;
		X1837 <= X1837;
		X1838 <= X1838;
		X1839 <= X1839;
		X1840 <= X1840;
		X1841 <= X1841;
		X1842 <= X1842;
		X1843 <= X1843;
		X1844 <= X1844;
		X1845 <= X1845;
		X1846 <= X1846;
		X1847 <= X1847;
		X1848 <= X1848;
		X1849 <= X1849;
		X1850 <= X1850;
		X1851 <= X1851;
		X1852 <= X1852;
		X1853 <= X1853;
		X1854 <= X1854;
		X1855 <= X1855;
		X1856 <= X1856;
		X1857 <= X1857;
		X1858 <= X1858;
		X1859 <= X1859;
		X1860 <= X1860;
		X1861 <= X1861;
		X1862 <= X1862;
		X1863 <= X1863;
		X1864 <= X1864;
		X1865 <= X1865;
		X1866 <= X1866;
		X1867 <= X1867;
		X1868 <= X1868;
		X1869 <= X1869;
		X1870 <= X1870;
		X1871 <= X1871;
		X1872 <= X1872;
		X1873 <= X1873;
		X1874 <= X1874;
		X1875 <= X1875;
		X1876 <= X1876;
		X1877 <= X1877;
		X1878 <= X1878;
		X1879 <= X1879;
		X1880 <= X1880;
		X1881 <= X1881;
		X1882 <= X1882;
		X1883 <= X1883;
		X1884 <= X1884;
		X1885 <= X1885;
		X1886 <= X1886;
		X1887 <= X1887;
		X1888 <= X1888;
		X1889 <= X1889;
		X1890 <= X1890;
		X1891 <= X1891;
		X1892 <= X1892;
		X1893 <= X1893;
		X1894 <= X1894;
		X1895 <= X1895;
		X1896 <= X1896;
		X1897 <= X1897;
		X1898 <= X1898;
		X1899 <= X1899;
		X1900 <= X1900;
		X1901 <= X1901;
		X1902 <= X1902;
		X1903 <= X1903;
		X1904 <= X1904;
		X1905 <= X1905;
		X1906 <= X1906;
		X1907 <= X1907;
		X1908 <= X1908;
		X1909 <= X1909;
		X1910 <= X1910;
		X1911 <= X1911;
		X1912 <= X1912;
		X1913 <= X1913;
		X1914 <= X1914;
		X1915 <= X1915;
		X1916 <= X1916;
		X1917 <= X1917;
		X1918 <= X1918;
		X1919 <= X1919;
		X1920 <= X1920;
		X1921 <= X1921;
		X1922 <= X1922;
		X1923 <= X1923;
		X1924 <= X1924;
		X1925 <= X1925;
		X1926 <= X1926;
		X1927 <= X1927;
		X1928 <= X1928;
		X1929 <= X1929;
		X1930 <= X1930;
		X1931 <= X1931;
		X1932 <= X1932;
		X1933 <= X1933;
		X1934 <= X1934;
		X1935 <= X1935;
		X1936 <= X1936;
		X1937 <= X1937;
		X1938 <= X1938;
		X1939 <= X1939;
		X1940 <= X1940;
		X1941 <= X1941;
		X1942 <= X1942;
		X1943 <= X1943;
		X1944 <= X1944;
		X1945 <= X1945;
		X1946 <= X1946;
		X1947 <= X1947;
		X1948 <= X1948;
		X1949 <= X1949;
		X1950 <= X1950;
		X1951 <= X1951;
		X1952 <= X1952;
		X1953 <= X1953;
		X1954 <= X1954;
		X1955 <= X1955;
		X1956 <= X1956;
		X1957 <= X1957;
		X1958 <= X1958;
		X1959 <= X1959;
		X1960 <= X1960;
		X1961 <= X1961;
		X1962 <= X1962;
		X1963 <= X1963;
		X1964 <= X1964;
		X1965 <= X1965;
		X1966 <= X1966;
		X1967 <= X1967;
		X1968 <= X1968;
		X1969 <= X1969;
		X1970 <= X1970;
		X1971 <= X1971;
		X1972 <= X1972;
		X1973 <= X1973;
		X1974 <= X1974;
		X1975 <= X1975;
		X1976 <= X1976;
		X1977 <= X1977;
		X1978 <= X1978;
		X1979 <= X1979;
		X1980 <= X1980;
		X1981 <= X1981;
		X1982 <= X1982;
		X1983 <= X1983;
		X1984 <= X1984;
		X1985 <= X1985;
		X1986 <= X1986;
		X1987 <= X1987;
		X1988 <= X1988;
		X1989 <= X1989;
		X1990 <= X1990;
		X1991 <= X1991;
		X1992 <= X1992;
		X1993 <= X1993;
		X1994 <= X1994;
		X1995 <= X1995;
		X1996 <= X1996;
		X1997 <= X1997;
		X1998 <= X1998;
		X1999 <= X1999;
		X2000 <= X2000;
		X2001 <= X2001;
		X2002 <= X2002;
		X2003 <= X2003;
		X2004 <= X2004;
		X2005 <= X2005;
		X2006 <= X2006;
		X2007 <= X2007;
		X2008 <= X2008;
		X2009 <= X2009;
		X2010 <= X2010;
		X2011 <= X2011;
		X2012 <= X2012;
		X2013 <= X2013;
		X2014 <= X2014;
		X2015 <= X2015;
		X2016 <= X2016;
		X2017 <= X2017;
		X2018 <= X2018;
		X2019 <= X2019;
		X2020 <= X2020;
		X2021 <= X2021;
		X2022 <= X2022;
		X2023 <= X2023;
		X2024 <= X2024;
		X2025 <= X2025;
		X2026 <= X2026;
		X2027 <= X2027;
		X2028 <= X2028;
		X2029 <= X2029;
		X2030 <= X2030;
		X2031 <= X2031;
		X2032 <= X2032;
		X2033 <= X2033;
		X2034 <= X2034;
		X2035 <= X2035;
		X2036 <= X2036;
		X2037 <= X2037;
		X2038 <= X2038;
		X2039 <= X2039;
		X2040 <= X2040;
		X2041 <= X2041;
		X2042 <= X2042;
		X2043 <= X2043;
		X2044 <= X2044;
		X2045 <= X2045;
		X2046 <= X2046;
		X2047 <= X2047);
	
	clock_control0 : clock_control
	PORT MAP();
	
		-- start_shiftin <= 
END interconnect;
