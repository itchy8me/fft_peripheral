LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
--USE IEEE.STD_LOGIC_ARITH.ALL;


--Shifts in 8 samples for parallel data ouput N=8 big
ENTITY c_2048to16x128_shifter IS
	PORT(
			--X0 downto X2048 ports input from ADC	
		X0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X4 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X5 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X6 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X7 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X8 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X9 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X10 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X11 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X12 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X13 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X14 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X15 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X16 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X17 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X18 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X19 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X20 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X21 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X22 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X23 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X24 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X25 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X26 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X27 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X28 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X29 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X30 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X31 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X32 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X33 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X34 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X35 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X36 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X37 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X38 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X39 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X40 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X41 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X42 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X43 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X44 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X45 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X46 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X47 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X48 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X49 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X50 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X51 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X52 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X53 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X54 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X55 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X56 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X57 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X58 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X59 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X60 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X61 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X62 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X63 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X64 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X65 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X66 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X67 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X68 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X69 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X70 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X71 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X72 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X73 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X74 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X75 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X76 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X77 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X78 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X79 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X80 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X81 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X82 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X83 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X84 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X85 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X86 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X87 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X88 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X89 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X90 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X91 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X92 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X93 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X94 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X95 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X96 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X97 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X98 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X99 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X100 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X101 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X102 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X103 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X104 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X105 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X106 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X107 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X108 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X109 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X110 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X111 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X112 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X113 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X114 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X115 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X116 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X117 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X118 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X119 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X120 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X121 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X122 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X123 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X124 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X125 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X126 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X127 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X128 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X129 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X130 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X131 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X132 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X133 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X134 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X135 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X136 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X137 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X138 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X139 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X140 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X141 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X142 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X143 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X144 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X145 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X146 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X147 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X148 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X149 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X150 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X151 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X152 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X153 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X154 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X155 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X156 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X157 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X158 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X159 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X160 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X161 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X162 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X163 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X164 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X165 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X166 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X167 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X168 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X169 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X170 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X171 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X172 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X173 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X174 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X175 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X176 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X177 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X178 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X179 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X180 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X181 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X182 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X183 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X184 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X185 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X186 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X187 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X188 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X189 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X190 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X191 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X192 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X193 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X194 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X195 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X196 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X197 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X198 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X199 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X200 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X201 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X202 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X203 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X204 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X205 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X206 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X207 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X208 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X209 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X210 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X211 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X212 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X213 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X214 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X215 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X216 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X217 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X218 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X219 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X220 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X221 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X222 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X223 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X224 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X225 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X226 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X227 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X228 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X229 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X230 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X231 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X232 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X233 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X234 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X235 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X236 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X237 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X238 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X239 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X240 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X241 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X242 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X243 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X244 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X245 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X246 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X247 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X248 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X249 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X250 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X251 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X252 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X253 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X254 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X255 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X256 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X257 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X258 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X259 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X260 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X261 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X262 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X263 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X264 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X265 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X266 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X267 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X268 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X269 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X270 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X271 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X272 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X273 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X274 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X275 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X276 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X277 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X278 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X279 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X280 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X281 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X282 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X283 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X284 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X285 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X286 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X287 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X288 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X289 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X290 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X291 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X292 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X293 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X294 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X295 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X296 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X297 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X298 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X299 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X300 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X301 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X302 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X303 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X304 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X305 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X306 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X307 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X308 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X309 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X310 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X311 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X312 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X313 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X314 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X315 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X316 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X317 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X318 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X319 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X320 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X321 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X322 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X323 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X324 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X325 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X326 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X327 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X328 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X329 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X330 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X331 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X332 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X333 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X334 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X335 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X336 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X337 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X338 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X339 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X340 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X341 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X342 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X343 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X344 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X345 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X346 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X347 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X348 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X349 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X350 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X351 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X352 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X353 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X354 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X355 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X356 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X357 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X358 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X359 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X360 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X361 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X362 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X363 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X364 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X365 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X366 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X367 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X368 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X369 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X370 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X371 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X372 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X373 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X374 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X375 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X376 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X377 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X378 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X379 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X380 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X381 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X382 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X383 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X384 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X385 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X386 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X387 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X388 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X389 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X390 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X391 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X392 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X393 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X394 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X395 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X396 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X397 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X398 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X399 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X400 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X401 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X402 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X403 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X404 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X405 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X406 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X407 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X408 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X409 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X410 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X411 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X412 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X413 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X414 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X415 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X416 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X417 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X418 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X419 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X420 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X421 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X422 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X423 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X424 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X425 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X426 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X427 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X428 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X429 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X430 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X431 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X432 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X433 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X434 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X435 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X436 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X437 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X438 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X439 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X440 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X441 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X442 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X443 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X444 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X445 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X446 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X447 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X448 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X449 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X450 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X451 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X452 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X453 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X454 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X455 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X456 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X457 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X458 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X459 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X460 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X461 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X462 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X463 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X464 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X465 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X466 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X467 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X468 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X469 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X470 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X471 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X472 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X473 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X474 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X475 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X476 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X477 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X478 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X479 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X480 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X481 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X482 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X483 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X484 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X485 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X486 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X487 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X488 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X489 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X490 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X491 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X492 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X493 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X494 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X495 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X496 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X497 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X498 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X499 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X500 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X501 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X502 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X503 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X504 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X505 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X506 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X507 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X508 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X509 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X510 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X511 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X512 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X513 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X514 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X515 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X516 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X517 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X518 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X519 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X520 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X521 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X522 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X523 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X524 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X525 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X526 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X527 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X528 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X529 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X530 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X531 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X532 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X533 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X534 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X535 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X536 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X537 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X538 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X539 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X540 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X541 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X542 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X543 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X544 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X545 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X546 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X547 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X548 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X549 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X550 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X551 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X552 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X553 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X554 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X555 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X556 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X557 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X558 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X559 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X560 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X561 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X562 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X563 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X564 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X565 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X566 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X567 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X568 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X569 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X570 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X571 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X572 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X573 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X574 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X575 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X576 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X577 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X578 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X579 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X580 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X581 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X582 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X583 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X584 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X585 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X586 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X587 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X588 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X589 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X590 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X591 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X592 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X593 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X594 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X595 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X596 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X597 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X598 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X599 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X600 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X601 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X602 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X603 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X604 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X605 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X606 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X607 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X608 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X609 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X610 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X611 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X612 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X613 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X614 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X615 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X616 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X617 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X618 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X619 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X620 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X621 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X622 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X623 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X624 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X625 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X626 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X627 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X628 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X629 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X630 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X631 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X632 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X633 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X634 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X635 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X636 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X637 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X638 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X639 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X640 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X641 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X642 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X643 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X644 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X645 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X646 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X647 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X648 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X649 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X650 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X651 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X652 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X653 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X654 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X655 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X656 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X657 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X658 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X659 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X660 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X661 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X662 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X663 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X664 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X665 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X666 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X667 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X668 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X669 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X670 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X671 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X672 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X673 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X674 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X675 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X676 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X677 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X678 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X679 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X680 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X681 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X682 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X683 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X684 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X685 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X686 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X687 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X688 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X689 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X690 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X691 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X692 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X693 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X694 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X695 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X696 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X697 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X698 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X699 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X700 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X701 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X702 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X703 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X704 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X705 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X706 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X707 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X708 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X709 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X710 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X711 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X712 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X713 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X714 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X715 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X716 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X717 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X718 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X719 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X720 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X721 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X722 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X723 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X724 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X725 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X726 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X727 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X728 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X729 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X730 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X731 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X732 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X733 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X734 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X735 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X736 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X737 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X738 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X739 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X740 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X741 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X742 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X743 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X744 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X745 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X746 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X747 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X748 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X749 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X750 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X751 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X752 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X753 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X754 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X755 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X756 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X757 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X758 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X759 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X760 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X761 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X762 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X763 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X764 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X765 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X766 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X767 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X768 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X769 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X770 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X771 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X772 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X773 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X774 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X775 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X776 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X777 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X778 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X779 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X780 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X781 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X782 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X783 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X784 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X785 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X786 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X787 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X788 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X789 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X790 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X791 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X792 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X793 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X794 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X795 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X796 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X797 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X798 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X799 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X800 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X801 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X802 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X803 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X804 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X805 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X806 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X807 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X808 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X809 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X810 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X811 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X812 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X813 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X814 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X815 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X816 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X817 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X818 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X819 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X820 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X821 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X822 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X823 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X824 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X825 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X826 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X827 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X828 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X829 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X830 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X831 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X832 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X833 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X834 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X835 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X836 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X837 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X838 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X839 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X840 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X841 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X842 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X843 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X844 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X845 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X846 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X847 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X848 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X849 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X850 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X851 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X852 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X853 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X854 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X855 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X856 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X857 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X858 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X859 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X860 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X861 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X862 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X863 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X864 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X865 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X866 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X867 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X868 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X869 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X870 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X871 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X872 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X873 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X874 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X875 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X876 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X877 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X878 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X879 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X880 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X881 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X882 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X883 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X884 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X885 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X886 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X887 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X888 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X889 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X890 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X891 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X892 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X893 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X894 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X895 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X896 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X897 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X898 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X899 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X900 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X901 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X902 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X903 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X904 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X905 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X906 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X907 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X908 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X909 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X910 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X911 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X912 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X913 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X914 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X915 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X916 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X917 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X918 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X919 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X920 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X921 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X922 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X923 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X924 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X925 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X926 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X927 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X928 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X929 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X930 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X931 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X932 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X933 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X934 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X935 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X936 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X937 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X938 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X939 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X940 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X941 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X942 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X943 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X944 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X945 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X946 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X947 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X948 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X949 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X950 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X951 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X952 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X953 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X954 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X955 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X956 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X957 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X958 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X959 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X960 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X961 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X962 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X963 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X964 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X965 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X966 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X967 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X968 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X969 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X970 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X971 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X972 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X973 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X974 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X975 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X976 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X977 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X978 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X979 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X980 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X981 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X982 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X983 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X984 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X985 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X986 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X987 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X988 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X989 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X990 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X991 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X992 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X993 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X994 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X995 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X996 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X997 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X998 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X999 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1000 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1001 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1002 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1003 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1004 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1005 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1006 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1007 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1008 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1009 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1010 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1011 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1012 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1013 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1014 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1015 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1016 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1017 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1018 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1019 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1020 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1021 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1022 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1023 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1024 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1025 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1026 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1027 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1028 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1029 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1030 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1031 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1032 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1033 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1034 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1035 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1036 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1037 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1038 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1039 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1040 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1041 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1042 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1043 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1044 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1045 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1046 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1047 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1048 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1049 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1050 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1051 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1052 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1053 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1054 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1055 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1056 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1057 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1058 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1059 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1060 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1061 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1062 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1063 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1064 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1065 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1066 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1067 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1068 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1069 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1070 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1071 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1072 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1073 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1074 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1075 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1076 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1077 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1078 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1079 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1080 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1081 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1082 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1083 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1084 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1085 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1086 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1087 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1088 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1089 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1090 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1091 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1092 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1093 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1094 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1095 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1096 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1097 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1098 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1099 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1100 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1101 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1102 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1103 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1104 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1105 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1106 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1107 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1108 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1109 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1110 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1111 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1112 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1113 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1114 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1115 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1116 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1117 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1118 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1119 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1120 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1121 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1122 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1123 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1124 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1125 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1126 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1127 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1128 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1129 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1130 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1131 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1132 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1133 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1134 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1135 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1136 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1137 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1138 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1139 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1140 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1141 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1142 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1143 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1144 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1145 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1146 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1147 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1148 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1149 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1150 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1151 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1152 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1153 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1154 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1155 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1156 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1157 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1158 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1159 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1160 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1161 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1162 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1163 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1164 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1165 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1166 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1167 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1168 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1169 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1170 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1171 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1172 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1173 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1174 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1175 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1176 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1177 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1178 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1179 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1180 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1181 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1182 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1183 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1184 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1185 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1186 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1187 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1188 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1189 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1190 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1191 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1192 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1193 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1194 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1195 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1196 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1197 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1198 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1199 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1200 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1201 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1202 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1203 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1204 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1205 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1206 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1207 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1208 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1209 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1210 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1211 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1212 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1213 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1214 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1215 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1216 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1217 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1218 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1219 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1220 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1221 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1222 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1223 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1224 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1225 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1226 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1227 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1228 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1229 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1230 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1231 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1232 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1233 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1234 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1235 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1236 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1237 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1238 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1239 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1240 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1241 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1242 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1243 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1244 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1245 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1246 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1247 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1248 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1249 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1250 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1251 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1252 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1253 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1254 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1255 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1256 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1257 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1258 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1259 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1260 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1261 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1262 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1263 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1264 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1265 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1266 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1267 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1268 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1269 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1270 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1271 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1272 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1273 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1274 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1275 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1276 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1277 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1278 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1279 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1280 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1281 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1282 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1283 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1284 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1285 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1286 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1287 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1288 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1289 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1290 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1291 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1292 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1293 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1294 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1295 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1296 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1297 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1298 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1299 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1300 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1301 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1302 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1303 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1304 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1305 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1306 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1307 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1308 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1309 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1310 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1311 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1312 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1313 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1314 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1315 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1316 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1317 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1318 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1319 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1320 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1321 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1322 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1323 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1324 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1325 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1326 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1327 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1328 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1329 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1330 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1331 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1332 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1333 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1334 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1335 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1336 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1337 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1338 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1339 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1340 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1341 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1342 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1343 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1344 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1345 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1346 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1347 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1348 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1349 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1350 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1351 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1352 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1353 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1354 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1355 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1356 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1357 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1358 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1359 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1360 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1361 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1362 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1363 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1364 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1365 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1366 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1367 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1368 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1369 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1370 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1371 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1372 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1373 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1374 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1375 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1376 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1377 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1378 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1379 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1380 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1381 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1382 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1383 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1384 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1385 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1386 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1387 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1388 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1389 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1390 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1391 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1392 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1393 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1394 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1395 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1396 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1397 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1398 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1399 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1400 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1401 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1402 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1403 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1404 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1405 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1406 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1407 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1408 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1409 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1410 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1411 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1412 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1413 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1414 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1415 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1416 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1417 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1418 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1419 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1420 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1421 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1422 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1423 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1424 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1425 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1426 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1427 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1428 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1429 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1430 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1431 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1432 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1433 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1434 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1435 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1436 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1437 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1438 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1439 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1440 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1441 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1442 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1443 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1444 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1445 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1446 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1447 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1448 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1449 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1450 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1451 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1452 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1453 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1454 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1455 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1456 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1457 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1458 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1459 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1460 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1461 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1462 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1463 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1464 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1465 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1466 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1467 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1468 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1469 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1470 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1471 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1472 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1473 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1474 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1475 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1476 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1477 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1478 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1479 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1480 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1481 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1482 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1483 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1484 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1485 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1486 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1487 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1488 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1489 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1490 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1491 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1492 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1493 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1494 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1495 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1496 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1497 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1498 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1499 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1500 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1501 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1502 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1503 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1504 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1505 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1506 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1507 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1508 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1509 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1510 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1511 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1512 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1513 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1514 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1515 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1516 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1517 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1518 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1519 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1520 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1521 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1522 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1523 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1524 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1525 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1526 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1527 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1528 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1529 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1530 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1531 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1532 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1533 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1534 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1535 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1536 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1537 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1538 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1539 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1540 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1541 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1542 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1543 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1544 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1545 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1546 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1547 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1548 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1549 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1550 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1551 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1552 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1553 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1554 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1555 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1556 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1557 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1558 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1559 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1560 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1561 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1562 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1563 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1564 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1565 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1566 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1567 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1568 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1569 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1570 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1571 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1572 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1573 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1574 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1575 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1576 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1577 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1578 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1579 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1580 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1581 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1582 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1583 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1584 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1585 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1586 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1587 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1588 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1589 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1590 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1591 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1592 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1593 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1594 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1595 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1596 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1597 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1598 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1599 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1600 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1601 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1602 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1603 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1604 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1605 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1606 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1607 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1608 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1609 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1610 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1611 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1612 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1613 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1614 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1615 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1616 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1617 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1618 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1619 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1620 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1621 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1622 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1623 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1624 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1625 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1626 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1627 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1628 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1629 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1630 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1631 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1632 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1633 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1634 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1635 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1636 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1637 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1638 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1639 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1640 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1641 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1642 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1643 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1644 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1645 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1646 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1647 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1648 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1649 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1650 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1651 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1652 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1653 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1654 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1655 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1656 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1657 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1658 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1659 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1660 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1661 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1662 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1663 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1664 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1665 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1666 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1667 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1668 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1669 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1670 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1671 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1672 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1673 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1674 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1675 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1676 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1677 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1678 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1679 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1680 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1681 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1682 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1683 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1684 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1685 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1686 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1687 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1688 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1689 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1690 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1691 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1692 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1693 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1694 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1695 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1696 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1697 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1698 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1699 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1700 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1701 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1702 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1703 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1704 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1705 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1706 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1707 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1708 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1709 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1710 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1711 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1712 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1713 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1714 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1715 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1716 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1717 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1718 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1719 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1720 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1721 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1722 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1723 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1724 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1725 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1726 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1727 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1728 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1729 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1730 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1731 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1732 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1733 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1734 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1735 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1736 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1737 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1738 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1739 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1740 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1741 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1742 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1743 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1744 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1745 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1746 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1747 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1748 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1749 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1750 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1751 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1752 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1753 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1754 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1755 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1756 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1757 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1758 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1759 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1760 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1761 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1762 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1763 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1764 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1765 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1766 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1767 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1768 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1769 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1770 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1771 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1772 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1773 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1774 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1775 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1776 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1777 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1778 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1779 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1780 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1781 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1782 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1783 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1784 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1785 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1786 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1787 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1788 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1789 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1790 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1791 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1792 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1793 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1794 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1795 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1796 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1797 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1798 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1799 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1800 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1801 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1802 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1803 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1804 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1805 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1806 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1807 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1808 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1809 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1810 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1811 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1812 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1813 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1814 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1815 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1816 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1817 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1818 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1819 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1820 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1821 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1822 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1823 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1824 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1825 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1826 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1827 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1828 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1829 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1830 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1831 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1832 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1833 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1834 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1835 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1836 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1837 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1838 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1839 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1840 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1841 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1842 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1843 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1844 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1845 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1846 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1847 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1848 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1849 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1850 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1851 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1852 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1853 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1854 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1855 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1856 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1857 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1858 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1859 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1860 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1861 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1862 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1863 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1864 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1865 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1866 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1867 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1868 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1869 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1870 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1871 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1872 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1873 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1874 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1875 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1876 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1877 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1878 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1879 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1880 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1881 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1882 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1883 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1884 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1885 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1886 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1887 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1888 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1889 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1890 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1891 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1892 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1893 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1894 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1895 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1896 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1897 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1898 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1899 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1900 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1901 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1902 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1903 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1904 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1905 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1906 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1907 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1908 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1909 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1910 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1911 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1912 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1913 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1914 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1915 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1916 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1917 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1918 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1919 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1920 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1921 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1922 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1923 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1924 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1925 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1926 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1927 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1928 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1929 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1930 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1931 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1932 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1933 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1934 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1935 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1936 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1937 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1938 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1939 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1940 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1941 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1942 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1943 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1944 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1945 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1946 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1947 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1948 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1949 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1950 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1951 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1952 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1953 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1954 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1955 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1956 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1957 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1958 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1959 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1960 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1961 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1962 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1963 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1964 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1965 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1966 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1967 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1968 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1969 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1970 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1971 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1972 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1973 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1974 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1975 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1976 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1977 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1978 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1979 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1980 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1981 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1982 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1983 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1984 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1985 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1986 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1987 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1988 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1989 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1990 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1991 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1992 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1993 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1994 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1995 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1996 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1997 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1998 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X1999 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2000 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2001 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2002 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2003 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2004 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2005 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2006 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2007 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2008 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2009 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2010 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2011 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2012 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2013 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2014 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2015 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2016 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2017 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2018 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2019 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2020 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2021 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2022 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2023 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2024 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2025 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2026 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2027 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2028 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2029 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2030 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2031 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2032 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2033 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2034 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2035 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2036 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2037 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2038 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2039 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2040 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2041 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2042 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2043 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2044 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2045 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2046 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		X2047 : IN STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		
		-- enable : IN STD_LOGIC := '0';
		FFT_finished : IN STD_LOGIC := '0';
		samples_ready : IN STD_LOGIC := '0';
		clk : IN STD_LOGIC := '0';
		
		-- sig_next : OUT STD_LOGIC := '0';
		shift_out0 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out1 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out2 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out3 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out4 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out5 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out6 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out7 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out8 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out9 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out10 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out11 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out12 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out13 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out14 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
		shift_out15 : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000");
END c_2048to16x128_shifter;


--the 4 bit to 7 bit (hex representation) decoding
ARCHITECTURE shift OF c_2048to16x128_shifter IS
	SIGNAL i : INTEGER := 0;
	-- SIGNAL data_incoming : STD_LOGIC := '0';
	
	SIGNAL XSIG0 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X0;
	SIGNAL XSIG1 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1;
	SIGNAL XSIG2 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2;
	SIGNAL XSIG3 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X3;
	SIGNAL XSIG4 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X4;
	SIGNAL XSIG5 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X5;
	SIGNAL XSIG6 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X6;
	SIGNAL XSIG7 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X7;
	SIGNAL XSIG8 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X8;
	SIGNAL XSIG9 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X9;
	SIGNAL XSIG10 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X10;
	SIGNAL XSIG11 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X11;
	SIGNAL XSIG12 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X12;
	SIGNAL XSIG13 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X13;
	SIGNAL XSIG14 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X14;
	SIGNAL XSIG15 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X15;
	SIGNAL XSIG16 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X16;
	SIGNAL XSIG17 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X17;
	SIGNAL XSIG18 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X18;
	SIGNAL XSIG19 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X19;
	SIGNAL XSIG20 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X20;
	SIGNAL XSIG21 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X21;
	SIGNAL XSIG22 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X22;
	SIGNAL XSIG23 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X23;
	SIGNAL XSIG24 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X24;
	SIGNAL XSIG25 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X25;
	SIGNAL XSIG26 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X26;
	SIGNAL XSIG27 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X27;
	SIGNAL XSIG28 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X28;
	SIGNAL XSIG29 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X29;
	SIGNAL XSIG30 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X30;
	SIGNAL XSIG31 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X31;
	SIGNAL XSIG32 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X32;
	SIGNAL XSIG33 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X33;
	SIGNAL XSIG34 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X34;
	SIGNAL XSIG35 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X35;
	SIGNAL XSIG36 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X36;
	SIGNAL XSIG37 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X37;
	SIGNAL XSIG38 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X38;
	SIGNAL XSIG39 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X39;
	SIGNAL XSIG40 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X40;
	SIGNAL XSIG41 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X41;
	SIGNAL XSIG42 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X42;
	SIGNAL XSIG43 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X43;
	SIGNAL XSIG44 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X44;
	SIGNAL XSIG45 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X45;
	SIGNAL XSIG46 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X46;
	SIGNAL XSIG47 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X47;
	SIGNAL XSIG48 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X48;
	SIGNAL XSIG49 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X49;
	SIGNAL XSIG50 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X50;
	SIGNAL XSIG51 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X51;
	SIGNAL XSIG52 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X52;
	SIGNAL XSIG53 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X53;
	SIGNAL XSIG54 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X54;
	SIGNAL XSIG55 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X55;
	SIGNAL XSIG56 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X56;
	SIGNAL XSIG57 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X57;
	SIGNAL XSIG58 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X58;
	SIGNAL XSIG59 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X59;
	SIGNAL XSIG60 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X60;
	SIGNAL XSIG61 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X61;
	SIGNAL XSIG62 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X62;
	SIGNAL XSIG63 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X63;
	SIGNAL XSIG64 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X64;
	SIGNAL XSIG65 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X65;
	SIGNAL XSIG66 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X66;
	SIGNAL XSIG67 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X67;
	SIGNAL XSIG68 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X68;
	SIGNAL XSIG69 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X69;
	SIGNAL XSIG70 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X70;
	SIGNAL XSIG71 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X71;
	SIGNAL XSIG72 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X72;
	SIGNAL XSIG73 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X73;
	SIGNAL XSIG74 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X74;
	SIGNAL XSIG75 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X75;
	SIGNAL XSIG76 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X76;
	SIGNAL XSIG77 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X77;
	SIGNAL XSIG78 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X78;
	SIGNAL XSIG79 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X79;
	SIGNAL XSIG80 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X80;
	SIGNAL XSIG81 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X81;
	SIGNAL XSIG82 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X82;
	SIGNAL XSIG83 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X83;
	SIGNAL XSIG84 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X84;
	SIGNAL XSIG85 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X85;
	SIGNAL XSIG86 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X86;
	SIGNAL XSIG87 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X87;
	SIGNAL XSIG88 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X88;
	SIGNAL XSIG89 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X89;
	SIGNAL XSIG90 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X90;
	SIGNAL XSIG91 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X91;
	SIGNAL XSIG92 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X92;
	SIGNAL XSIG93 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X93;
	SIGNAL XSIG94 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X94;
	SIGNAL XSIG95 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X95;
	SIGNAL XSIG96 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X96;
	SIGNAL XSIG97 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X97;
	SIGNAL XSIG98 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X98;
	SIGNAL XSIG99 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X99;
	SIGNAL XSIG100 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X100;
	SIGNAL XSIG101 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X101;
	SIGNAL XSIG102 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X102;
	SIGNAL XSIG103 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X103;
	SIGNAL XSIG104 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X104;
	SIGNAL XSIG105 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X105;
	SIGNAL XSIG106 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X106;
	SIGNAL XSIG107 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X107;
	SIGNAL XSIG108 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X108;
	SIGNAL XSIG109 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X109;
	SIGNAL XSIG110 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X110;
	SIGNAL XSIG111 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X111;
	SIGNAL XSIG112 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X112;
	SIGNAL XSIG113 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X113;
	SIGNAL XSIG114 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X114;
	SIGNAL XSIG115 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X115;
	SIGNAL XSIG116 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X116;
	SIGNAL XSIG117 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X117;
	SIGNAL XSIG118 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X118;
	SIGNAL XSIG119 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X119;
	SIGNAL XSIG120 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X120;
	SIGNAL XSIG121 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X121;
	SIGNAL XSIG122 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X122;
	SIGNAL XSIG123 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X123;
	SIGNAL XSIG124 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X124;
	SIGNAL XSIG125 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X125;
	SIGNAL XSIG126 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X126;
	SIGNAL XSIG127 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X127;
	SIGNAL XSIG128 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X128;
	SIGNAL XSIG129 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X129;
	SIGNAL XSIG130 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X130;
	SIGNAL XSIG131 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X131;
	SIGNAL XSIG132 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X132;
	SIGNAL XSIG133 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X133;
	SIGNAL XSIG134 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X134;
	SIGNAL XSIG135 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X135;
	SIGNAL XSIG136 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X136;
	SIGNAL XSIG137 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X137;
	SIGNAL XSIG138 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X138;
	SIGNAL XSIG139 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X139;
	SIGNAL XSIG140 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X140;
	SIGNAL XSIG141 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X141;
	SIGNAL XSIG142 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X142;
	SIGNAL XSIG143 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X143;
	SIGNAL XSIG144 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X144;
	SIGNAL XSIG145 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X145;
	SIGNAL XSIG146 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X146;
	SIGNAL XSIG147 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X147;
	SIGNAL XSIG148 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X148;
	SIGNAL XSIG149 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X149;
	SIGNAL XSIG150 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X150;
	SIGNAL XSIG151 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X151;
	SIGNAL XSIG152 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X152;
	SIGNAL XSIG153 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X153;
	SIGNAL XSIG154 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X154;
	SIGNAL XSIG155 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X155;
	SIGNAL XSIG156 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X156;
	SIGNAL XSIG157 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X157;
	SIGNAL XSIG158 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X158;
	SIGNAL XSIG159 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X159;
	SIGNAL XSIG160 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X160;
	SIGNAL XSIG161 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X161;
	SIGNAL XSIG162 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X162;
	SIGNAL XSIG163 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X163;
	SIGNAL XSIG164 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X164;
	SIGNAL XSIG165 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X165;
	SIGNAL XSIG166 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X166;
	SIGNAL XSIG167 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X167;
	SIGNAL XSIG168 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X168;
	SIGNAL XSIG169 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X169;
	SIGNAL XSIG170 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X170;
	SIGNAL XSIG171 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X171;
	SIGNAL XSIG172 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X172;
	SIGNAL XSIG173 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X173;
	SIGNAL XSIG174 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X174;
	SIGNAL XSIG175 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X175;
	SIGNAL XSIG176 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X176;
	SIGNAL XSIG177 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X177;
	SIGNAL XSIG178 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X178;
	SIGNAL XSIG179 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X179;
	SIGNAL XSIG180 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X180;
	SIGNAL XSIG181 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X181;
	SIGNAL XSIG182 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X182;
	SIGNAL XSIG183 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X183;
	SIGNAL XSIG184 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X184;
	SIGNAL XSIG185 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X185;
	SIGNAL XSIG186 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X186;
	SIGNAL XSIG187 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X187;
	SIGNAL XSIG188 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X188;
	SIGNAL XSIG189 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X189;
	SIGNAL XSIG190 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X190;
	SIGNAL XSIG191 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X191;
	SIGNAL XSIG192 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X192;
	SIGNAL XSIG193 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X193;
	SIGNAL XSIG194 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X194;
	SIGNAL XSIG195 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X195;
	SIGNAL XSIG196 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X196;
	SIGNAL XSIG197 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X197;
	SIGNAL XSIG198 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X198;
	SIGNAL XSIG199 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X199;
	SIGNAL XSIG200 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X200;
	SIGNAL XSIG201 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X201;
	SIGNAL XSIG202 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X202;
	SIGNAL XSIG203 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X203;
	SIGNAL XSIG204 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X204;
	SIGNAL XSIG205 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X205;
	SIGNAL XSIG206 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X206;
	SIGNAL XSIG207 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X207;
	SIGNAL XSIG208 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X208;
	SIGNAL XSIG209 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X209;
	SIGNAL XSIG210 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X210;
	SIGNAL XSIG211 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X211;
	SIGNAL XSIG212 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X212;
	SIGNAL XSIG213 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X213;
	SIGNAL XSIG214 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X214;
	SIGNAL XSIG215 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X215;
	SIGNAL XSIG216 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X216;
	SIGNAL XSIG217 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X217;
	SIGNAL XSIG218 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X218;
	SIGNAL XSIG219 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X219;
	SIGNAL XSIG220 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X220;
	SIGNAL XSIG221 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X221;
	SIGNAL XSIG222 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X222;
	SIGNAL XSIG223 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X223;
	SIGNAL XSIG224 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X224;
	SIGNAL XSIG225 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X225;
	SIGNAL XSIG226 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X226;
	SIGNAL XSIG227 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X227;
	SIGNAL XSIG228 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X228;
	SIGNAL XSIG229 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X229;
	SIGNAL XSIG230 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X230;
	SIGNAL XSIG231 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X231;
	SIGNAL XSIG232 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X232;
	SIGNAL XSIG233 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X233;
	SIGNAL XSIG234 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X234;
	SIGNAL XSIG235 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X235;
	SIGNAL XSIG236 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X236;
	SIGNAL XSIG237 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X237;
	SIGNAL XSIG238 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X238;
	SIGNAL XSIG239 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X239;
	SIGNAL XSIG240 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X240;
	SIGNAL XSIG241 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X241;
	SIGNAL XSIG242 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X242;
	SIGNAL XSIG243 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X243;
	SIGNAL XSIG244 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X244;
	SIGNAL XSIG245 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X245;
	SIGNAL XSIG246 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X246;
	SIGNAL XSIG247 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X247;
	SIGNAL XSIG248 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X248;
	SIGNAL XSIG249 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X249;
	SIGNAL XSIG250 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X250;
	SIGNAL XSIG251 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X251;
	SIGNAL XSIG252 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X252;
	SIGNAL XSIG253 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X253;
	SIGNAL XSIG254 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X254;
	SIGNAL XSIG255 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X255;
	SIGNAL XSIG256 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X256;
	SIGNAL XSIG257 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X257;
	SIGNAL XSIG258 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X258;
	SIGNAL XSIG259 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X259;
	SIGNAL XSIG260 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X260;
	SIGNAL XSIG261 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X261;
	SIGNAL XSIG262 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X262;
	SIGNAL XSIG263 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X263;
	SIGNAL XSIG264 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X264;
	SIGNAL XSIG265 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X265;
	SIGNAL XSIG266 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X266;
	SIGNAL XSIG267 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X267;
	SIGNAL XSIG268 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X268;
	SIGNAL XSIG269 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X269;
	SIGNAL XSIG270 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X270;
	SIGNAL XSIG271 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X271;
	SIGNAL XSIG272 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X272;
	SIGNAL XSIG273 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X273;
	SIGNAL XSIG274 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X274;
	SIGNAL XSIG275 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X275;
	SIGNAL XSIG276 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X276;
	SIGNAL XSIG277 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X277;
	SIGNAL XSIG278 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X278;
	SIGNAL XSIG279 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X279;
	SIGNAL XSIG280 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X280;
	SIGNAL XSIG281 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X281;
	SIGNAL XSIG282 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X282;
	SIGNAL XSIG283 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X283;
	SIGNAL XSIG284 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X284;
	SIGNAL XSIG285 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X285;
	SIGNAL XSIG286 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X286;
	SIGNAL XSIG287 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X287;
	SIGNAL XSIG288 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X288;
	SIGNAL XSIG289 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X289;
	SIGNAL XSIG290 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X290;
	SIGNAL XSIG291 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X291;
	SIGNAL XSIG292 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X292;
	SIGNAL XSIG293 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X293;
	SIGNAL XSIG294 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X294;
	SIGNAL XSIG295 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X295;
	SIGNAL XSIG296 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X296;
	SIGNAL XSIG297 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X297;
	SIGNAL XSIG298 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X298;
	SIGNAL XSIG299 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X299;
	SIGNAL XSIG300 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X300;
	SIGNAL XSIG301 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X301;
	SIGNAL XSIG302 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X302;
	SIGNAL XSIG303 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X303;
	SIGNAL XSIG304 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X304;
	SIGNAL XSIG305 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X305;
	SIGNAL XSIG306 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X306;
	SIGNAL XSIG307 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X307;
	SIGNAL XSIG308 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X308;
	SIGNAL XSIG309 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X309;
	SIGNAL XSIG310 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X310;
	SIGNAL XSIG311 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X311;
	SIGNAL XSIG312 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X312;
	SIGNAL XSIG313 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X313;
	SIGNAL XSIG314 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X314;
	SIGNAL XSIG315 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X315;
	SIGNAL XSIG316 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X316;
	SIGNAL XSIG317 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X317;
	SIGNAL XSIG318 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X318;
	SIGNAL XSIG319 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X319;
	SIGNAL XSIG320 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X320;
	SIGNAL XSIG321 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X321;
	SIGNAL XSIG322 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X322;
	SIGNAL XSIG323 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X323;
	SIGNAL XSIG324 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X324;
	SIGNAL XSIG325 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X325;
	SIGNAL XSIG326 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X326;
	SIGNAL XSIG327 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X327;
	SIGNAL XSIG328 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X328;
	SIGNAL XSIG329 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X329;
	SIGNAL XSIG330 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X330;
	SIGNAL XSIG331 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X331;
	SIGNAL XSIG332 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X332;
	SIGNAL XSIG333 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X333;
	SIGNAL XSIG334 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X334;
	SIGNAL XSIG335 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X335;
	SIGNAL XSIG336 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X336;
	SIGNAL XSIG337 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X337;
	SIGNAL XSIG338 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X338;
	SIGNAL XSIG339 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X339;
	SIGNAL XSIG340 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X340;
	SIGNAL XSIG341 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X341;
	SIGNAL XSIG342 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X342;
	SIGNAL XSIG343 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X343;
	SIGNAL XSIG344 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X344;
	SIGNAL XSIG345 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X345;
	SIGNAL XSIG346 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X346;
	SIGNAL XSIG347 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X347;
	SIGNAL XSIG348 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X348;
	SIGNAL XSIG349 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X349;
	SIGNAL XSIG350 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X350;
	SIGNAL XSIG351 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X351;
	SIGNAL XSIG352 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X352;
	SIGNAL XSIG353 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X353;
	SIGNAL XSIG354 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X354;
	SIGNAL XSIG355 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X355;
	SIGNAL XSIG356 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X356;
	SIGNAL XSIG357 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X357;
	SIGNAL XSIG358 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X358;
	SIGNAL XSIG359 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X359;
	SIGNAL XSIG360 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X360;
	SIGNAL XSIG361 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X361;
	SIGNAL XSIG362 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X362;
	SIGNAL XSIG363 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X363;
	SIGNAL XSIG364 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X364;
	SIGNAL XSIG365 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X365;
	SIGNAL XSIG366 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X366;
	SIGNAL XSIG367 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X367;
	SIGNAL XSIG368 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X368;
	SIGNAL XSIG369 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X369;
	SIGNAL XSIG370 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X370;
	SIGNAL XSIG371 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X371;
	SIGNAL XSIG372 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X372;
	SIGNAL XSIG373 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X373;
	SIGNAL XSIG374 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X374;
	SIGNAL XSIG375 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X375;
	SIGNAL XSIG376 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X376;
	SIGNAL XSIG377 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X377;
	SIGNAL XSIG378 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X378;
	SIGNAL XSIG379 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X379;
	SIGNAL XSIG380 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X380;
	SIGNAL XSIG381 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X381;
	SIGNAL XSIG382 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X382;
	SIGNAL XSIG383 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X383;
	SIGNAL XSIG384 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X384;
	SIGNAL XSIG385 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X385;
	SIGNAL XSIG386 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X386;
	SIGNAL XSIG387 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X387;
	SIGNAL XSIG388 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X388;
	SIGNAL XSIG389 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X389;
	SIGNAL XSIG390 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X390;
	SIGNAL XSIG391 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X391;
	SIGNAL XSIG392 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X392;
	SIGNAL XSIG393 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X393;
	SIGNAL XSIG394 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X394;
	SIGNAL XSIG395 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X395;
	SIGNAL XSIG396 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X396;
	SIGNAL XSIG397 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X397;
	SIGNAL XSIG398 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X398;
	SIGNAL XSIG399 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X399;
	SIGNAL XSIG400 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X400;
	SIGNAL XSIG401 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X401;
	SIGNAL XSIG402 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X402;
	SIGNAL XSIG403 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X403;
	SIGNAL XSIG404 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X404;
	SIGNAL XSIG405 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X405;
	SIGNAL XSIG406 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X406;
	SIGNAL XSIG407 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X407;
	SIGNAL XSIG408 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X408;
	SIGNAL XSIG409 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X409;
	SIGNAL XSIG410 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X410;
	SIGNAL XSIG411 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X411;
	SIGNAL XSIG412 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X412;
	SIGNAL XSIG413 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X413;
	SIGNAL XSIG414 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X414;
	SIGNAL XSIG415 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X415;
	SIGNAL XSIG416 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X416;
	SIGNAL XSIG417 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X417;
	SIGNAL XSIG418 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X418;
	SIGNAL XSIG419 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X419;
	SIGNAL XSIG420 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X420;
	SIGNAL XSIG421 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X421;
	SIGNAL XSIG422 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X422;
	SIGNAL XSIG423 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X423;
	SIGNAL XSIG424 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X424;
	SIGNAL XSIG425 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X425;
	SIGNAL XSIG426 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X426;
	SIGNAL XSIG427 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X427;
	SIGNAL XSIG428 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X428;
	SIGNAL XSIG429 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X429;
	SIGNAL XSIG430 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X430;
	SIGNAL XSIG431 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X431;
	SIGNAL XSIG432 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X432;
	SIGNAL XSIG433 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X433;
	SIGNAL XSIG434 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X434;
	SIGNAL XSIG435 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X435;
	SIGNAL XSIG436 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X436;
	SIGNAL XSIG437 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X437;
	SIGNAL XSIG438 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X438;
	SIGNAL XSIG439 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X439;
	SIGNAL XSIG440 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X440;
	SIGNAL XSIG441 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X441;
	SIGNAL XSIG442 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X442;
	SIGNAL XSIG443 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X443;
	SIGNAL XSIG444 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X444;
	SIGNAL XSIG445 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X445;
	SIGNAL XSIG446 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X446;
	SIGNAL XSIG447 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X447;
	SIGNAL XSIG448 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X448;
	SIGNAL XSIG449 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X449;
	SIGNAL XSIG450 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X450;
	SIGNAL XSIG451 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X451;
	SIGNAL XSIG452 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X452;
	SIGNAL XSIG453 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X453;
	SIGNAL XSIG454 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X454;
	SIGNAL XSIG455 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X455;
	SIGNAL XSIG456 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X456;
	SIGNAL XSIG457 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X457;
	SIGNAL XSIG458 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X458;
	SIGNAL XSIG459 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X459;
	SIGNAL XSIG460 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X460;
	SIGNAL XSIG461 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X461;
	SIGNAL XSIG462 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X462;
	SIGNAL XSIG463 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X463;
	SIGNAL XSIG464 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X464;
	SIGNAL XSIG465 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X465;
	SIGNAL XSIG466 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X466;
	SIGNAL XSIG467 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X467;
	SIGNAL XSIG468 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X468;
	SIGNAL XSIG469 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X469;
	SIGNAL XSIG470 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X470;
	SIGNAL XSIG471 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X471;
	SIGNAL XSIG472 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X472;
	SIGNAL XSIG473 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X473;
	SIGNAL XSIG474 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X474;
	SIGNAL XSIG475 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X475;
	SIGNAL XSIG476 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X476;
	SIGNAL XSIG477 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X477;
	SIGNAL XSIG478 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X478;
	SIGNAL XSIG479 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X479;
	SIGNAL XSIG480 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X480;
	SIGNAL XSIG481 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X481;
	SIGNAL XSIG482 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X482;
	SIGNAL XSIG483 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X483;
	SIGNAL XSIG484 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X484;
	SIGNAL XSIG485 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X485;
	SIGNAL XSIG486 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X486;
	SIGNAL XSIG487 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X487;
	SIGNAL XSIG488 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X488;
	SIGNAL XSIG489 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X489;
	SIGNAL XSIG490 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X490;
	SIGNAL XSIG491 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X491;
	SIGNAL XSIG492 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X492;
	SIGNAL XSIG493 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X493;
	SIGNAL XSIG494 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X494;
	SIGNAL XSIG495 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X495;
	SIGNAL XSIG496 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X496;
	SIGNAL XSIG497 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X497;
	SIGNAL XSIG498 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X498;
	SIGNAL XSIG499 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X499;
	SIGNAL XSIG500 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X500;
	SIGNAL XSIG501 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X501;
	SIGNAL XSIG502 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X502;
	SIGNAL XSIG503 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X503;
	SIGNAL XSIG504 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X504;
	SIGNAL XSIG505 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X505;
	SIGNAL XSIG506 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X506;
	SIGNAL XSIG507 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X507;
	SIGNAL XSIG508 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X508;
	SIGNAL XSIG509 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X509;
	SIGNAL XSIG510 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X510;
	SIGNAL XSIG511 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X511;
	SIGNAL XSIG512 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X512;
	SIGNAL XSIG513 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X513;
	SIGNAL XSIG514 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X514;
	SIGNAL XSIG515 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X515;
	SIGNAL XSIG516 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X516;
	SIGNAL XSIG517 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X517;
	SIGNAL XSIG518 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X518;
	SIGNAL XSIG519 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X519;
	SIGNAL XSIG520 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X520;
	SIGNAL XSIG521 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X521;
	SIGNAL XSIG522 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X522;
	SIGNAL XSIG523 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X523;
	SIGNAL XSIG524 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X524;
	SIGNAL XSIG525 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X525;
	SIGNAL XSIG526 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X526;
	SIGNAL XSIG527 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X527;
	SIGNAL XSIG528 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X528;
	SIGNAL XSIG529 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X529;
	SIGNAL XSIG530 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X530;
	SIGNAL XSIG531 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X531;
	SIGNAL XSIG532 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X532;
	SIGNAL XSIG533 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X533;
	SIGNAL XSIG534 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X534;
	SIGNAL XSIG535 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X535;
	SIGNAL XSIG536 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X536;
	SIGNAL XSIG537 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X537;
	SIGNAL XSIG538 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X538;
	SIGNAL XSIG539 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X539;
	SIGNAL XSIG540 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X540;
	SIGNAL XSIG541 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X541;
	SIGNAL XSIG542 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X542;
	SIGNAL XSIG543 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X543;
	SIGNAL XSIG544 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X544;
	SIGNAL XSIG545 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X545;
	SIGNAL XSIG546 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X546;
	SIGNAL XSIG547 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X547;
	SIGNAL XSIG548 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X548;
	SIGNAL XSIG549 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X549;
	SIGNAL XSIG550 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X550;
	SIGNAL XSIG551 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X551;
	SIGNAL XSIG552 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X552;
	SIGNAL XSIG553 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X553;
	SIGNAL XSIG554 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X554;
	SIGNAL XSIG555 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X555;
	SIGNAL XSIG556 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X556;
	SIGNAL XSIG557 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X557;
	SIGNAL XSIG558 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X558;
	SIGNAL XSIG559 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X559;
	SIGNAL XSIG560 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X560;
	SIGNAL XSIG561 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X561;
	SIGNAL XSIG562 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X562;
	SIGNAL XSIG563 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X563;
	SIGNAL XSIG564 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X564;
	SIGNAL XSIG565 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X565;
	SIGNAL XSIG566 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X566;
	SIGNAL XSIG567 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X567;
	SIGNAL XSIG568 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X568;
	SIGNAL XSIG569 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X569;
	SIGNAL XSIG570 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X570;
	SIGNAL XSIG571 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X571;
	SIGNAL XSIG572 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X572;
	SIGNAL XSIG573 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X573;
	SIGNAL XSIG574 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X574;
	SIGNAL XSIG575 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X575;
	SIGNAL XSIG576 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X576;
	SIGNAL XSIG577 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X577;
	SIGNAL XSIG578 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X578;
	SIGNAL XSIG579 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X579;
	SIGNAL XSIG580 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X580;
	SIGNAL XSIG581 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X581;
	SIGNAL XSIG582 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X582;
	SIGNAL XSIG583 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X583;
	SIGNAL XSIG584 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X584;
	SIGNAL XSIG585 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X585;
	SIGNAL XSIG586 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X586;
	SIGNAL XSIG587 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X587;
	SIGNAL XSIG588 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X588;
	SIGNAL XSIG589 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X589;
	SIGNAL XSIG590 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X590;
	SIGNAL XSIG591 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X591;
	SIGNAL XSIG592 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X592;
	SIGNAL XSIG593 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X593;
	SIGNAL XSIG594 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X594;
	SIGNAL XSIG595 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X595;
	SIGNAL XSIG596 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X596;
	SIGNAL XSIG597 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X597;
	SIGNAL XSIG598 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X598;
	SIGNAL XSIG599 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X599;
	SIGNAL XSIG600 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X600;
	SIGNAL XSIG601 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X601;
	SIGNAL XSIG602 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X602;
	SIGNAL XSIG603 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X603;
	SIGNAL XSIG604 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X604;
	SIGNAL XSIG605 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X605;
	SIGNAL XSIG606 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X606;
	SIGNAL XSIG607 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X607;
	SIGNAL XSIG608 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X608;
	SIGNAL XSIG609 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X609;
	SIGNAL XSIG610 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X610;
	SIGNAL XSIG611 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X611;
	SIGNAL XSIG612 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X612;
	SIGNAL XSIG613 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X613;
	SIGNAL XSIG614 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X614;
	SIGNAL XSIG615 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X615;
	SIGNAL XSIG616 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X616;
	SIGNAL XSIG617 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X617;
	SIGNAL XSIG618 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X618;
	SIGNAL XSIG619 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X619;
	SIGNAL XSIG620 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X620;
	SIGNAL XSIG621 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X621;
	SIGNAL XSIG622 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X622;
	SIGNAL XSIG623 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X623;
	SIGNAL XSIG624 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X624;
	SIGNAL XSIG625 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X625;
	SIGNAL XSIG626 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X626;
	SIGNAL XSIG627 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X627;
	SIGNAL XSIG628 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X628;
	SIGNAL XSIG629 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X629;
	SIGNAL XSIG630 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X630;
	SIGNAL XSIG631 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X631;
	SIGNAL XSIG632 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X632;
	SIGNAL XSIG633 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X633;
	SIGNAL XSIG634 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X634;
	SIGNAL XSIG635 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X635;
	SIGNAL XSIG636 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X636;
	SIGNAL XSIG637 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X637;
	SIGNAL XSIG638 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X638;
	SIGNAL XSIG639 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X639;
	SIGNAL XSIG640 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X640;
	SIGNAL XSIG641 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X641;
	SIGNAL XSIG642 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X642;
	SIGNAL XSIG643 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X643;
	SIGNAL XSIG644 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X644;
	SIGNAL XSIG645 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X645;
	SIGNAL XSIG646 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X646;
	SIGNAL XSIG647 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X647;
	SIGNAL XSIG648 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X648;
	SIGNAL XSIG649 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X649;
	SIGNAL XSIG650 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X650;
	SIGNAL XSIG651 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X651;
	SIGNAL XSIG652 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X652;
	SIGNAL XSIG653 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X653;
	SIGNAL XSIG654 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X654;
	SIGNAL XSIG655 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X655;
	SIGNAL XSIG656 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X656;
	SIGNAL XSIG657 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X657;
	SIGNAL XSIG658 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X658;
	SIGNAL XSIG659 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X659;
	SIGNAL XSIG660 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X660;
	SIGNAL XSIG661 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X661;
	SIGNAL XSIG662 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X662;
	SIGNAL XSIG663 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X663;
	SIGNAL XSIG664 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X664;
	SIGNAL XSIG665 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X665;
	SIGNAL XSIG666 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X666;
	SIGNAL XSIG667 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X667;
	SIGNAL XSIG668 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X668;
	SIGNAL XSIG669 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X669;
	SIGNAL XSIG670 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X670;
	SIGNAL XSIG671 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X671;
	SIGNAL XSIG672 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X672;
	SIGNAL XSIG673 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X673;
	SIGNAL XSIG674 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X674;
	SIGNAL XSIG675 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X675;
	SIGNAL XSIG676 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X676;
	SIGNAL XSIG677 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X677;
	SIGNAL XSIG678 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X678;
	SIGNAL XSIG679 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X679;
	SIGNAL XSIG680 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X680;
	SIGNAL XSIG681 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X681;
	SIGNAL XSIG682 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X682;
	SIGNAL XSIG683 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X683;
	SIGNAL XSIG684 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X684;
	SIGNAL XSIG685 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X685;
	SIGNAL XSIG686 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X686;
	SIGNAL XSIG687 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X687;
	SIGNAL XSIG688 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X688;
	SIGNAL XSIG689 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X689;
	SIGNAL XSIG690 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X690;
	SIGNAL XSIG691 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X691;
	SIGNAL XSIG692 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X692;
	SIGNAL XSIG693 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X693;
	SIGNAL XSIG694 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X694;
	SIGNAL XSIG695 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X695;
	SIGNAL XSIG696 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X696;
	SIGNAL XSIG697 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X697;
	SIGNAL XSIG698 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X698;
	SIGNAL XSIG699 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X699;
	SIGNAL XSIG700 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X700;
	SIGNAL XSIG701 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X701;
	SIGNAL XSIG702 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X702;
	SIGNAL XSIG703 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X703;
	SIGNAL XSIG704 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X704;
	SIGNAL XSIG705 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X705;
	SIGNAL XSIG706 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X706;
	SIGNAL XSIG707 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X707;
	SIGNAL XSIG708 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X708;
	SIGNAL XSIG709 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X709;
	SIGNAL XSIG710 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X710;
	SIGNAL XSIG711 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X711;
	SIGNAL XSIG712 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X712;
	SIGNAL XSIG713 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X713;
	SIGNAL XSIG714 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X714;
	SIGNAL XSIG715 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X715;
	SIGNAL XSIG716 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X716;
	SIGNAL XSIG717 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X717;
	SIGNAL XSIG718 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X718;
	SIGNAL XSIG719 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X719;
	SIGNAL XSIG720 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X720;
	SIGNAL XSIG721 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X721;
	SIGNAL XSIG722 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X722;
	SIGNAL XSIG723 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X723;
	SIGNAL XSIG724 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X724;
	SIGNAL XSIG725 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X725;
	SIGNAL XSIG726 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X726;
	SIGNAL XSIG727 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X727;
	SIGNAL XSIG728 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X728;
	SIGNAL XSIG729 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X729;
	SIGNAL XSIG730 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X730;
	SIGNAL XSIG731 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X731;
	SIGNAL XSIG732 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X732;
	SIGNAL XSIG733 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X733;
	SIGNAL XSIG734 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X734;
	SIGNAL XSIG735 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X735;
	SIGNAL XSIG736 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X736;
	SIGNAL XSIG737 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X737;
	SIGNAL XSIG738 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X738;
	SIGNAL XSIG739 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X739;
	SIGNAL XSIG740 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X740;
	SIGNAL XSIG741 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X741;
	SIGNAL XSIG742 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X742;
	SIGNAL XSIG743 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X743;
	SIGNAL XSIG744 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X744;
	SIGNAL XSIG745 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X745;
	SIGNAL XSIG746 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X746;
	SIGNAL XSIG747 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X747;
	SIGNAL XSIG748 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X748;
	SIGNAL XSIG749 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X749;
	SIGNAL XSIG750 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X750;
	SIGNAL XSIG751 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X751;
	SIGNAL XSIG752 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X752;
	SIGNAL XSIG753 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X753;
	SIGNAL XSIG754 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X754;
	SIGNAL XSIG755 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X755;
	SIGNAL XSIG756 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X756;
	SIGNAL XSIG757 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X757;
	SIGNAL XSIG758 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X758;
	SIGNAL XSIG759 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X759;
	SIGNAL XSIG760 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X760;
	SIGNAL XSIG761 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X761;
	SIGNAL XSIG762 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X762;
	SIGNAL XSIG763 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X763;
	SIGNAL XSIG764 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X764;
	SIGNAL XSIG765 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X765;
	SIGNAL XSIG766 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X766;
	SIGNAL XSIG767 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X767;
	SIGNAL XSIG768 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X768;
	SIGNAL XSIG769 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X769;
	SIGNAL XSIG770 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X770;
	SIGNAL XSIG771 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X771;
	SIGNAL XSIG772 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X772;
	SIGNAL XSIG773 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X773;
	SIGNAL XSIG774 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X774;
	SIGNAL XSIG775 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X775;
	SIGNAL XSIG776 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X776;
	SIGNAL XSIG777 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X777;
	SIGNAL XSIG778 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X778;
	SIGNAL XSIG779 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X779;
	SIGNAL XSIG780 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X780;
	SIGNAL XSIG781 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X781;
	SIGNAL XSIG782 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X782;
	SIGNAL XSIG783 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X783;
	SIGNAL XSIG784 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X784;
	SIGNAL XSIG785 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X785;
	SIGNAL XSIG786 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X786;
	SIGNAL XSIG787 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X787;
	SIGNAL XSIG788 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X788;
	SIGNAL XSIG789 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X789;
	SIGNAL XSIG790 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X790;
	SIGNAL XSIG791 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X791;
	SIGNAL XSIG792 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X792;
	SIGNAL XSIG793 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X793;
	SIGNAL XSIG794 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X794;
	SIGNAL XSIG795 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X795;
	SIGNAL XSIG796 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X796;
	SIGNAL XSIG797 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X797;
	SIGNAL XSIG798 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X798;
	SIGNAL XSIG799 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X799;
	SIGNAL XSIG800 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X800;
	SIGNAL XSIG801 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X801;
	SIGNAL XSIG802 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X802;
	SIGNAL XSIG803 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X803;
	SIGNAL XSIG804 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X804;
	SIGNAL XSIG805 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X805;
	SIGNAL XSIG806 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X806;
	SIGNAL XSIG807 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X807;
	SIGNAL XSIG808 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X808;
	SIGNAL XSIG809 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X809;
	SIGNAL XSIG810 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X810;
	SIGNAL XSIG811 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X811;
	SIGNAL XSIG812 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X812;
	SIGNAL XSIG813 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X813;
	SIGNAL XSIG814 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X814;
	SIGNAL XSIG815 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X815;
	SIGNAL XSIG816 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X816;
	SIGNAL XSIG817 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X817;
	SIGNAL XSIG818 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X818;
	SIGNAL XSIG819 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X819;
	SIGNAL XSIG820 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X820;
	SIGNAL XSIG821 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X821;
	SIGNAL XSIG822 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X822;
	SIGNAL XSIG823 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X823;
	SIGNAL XSIG824 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X824;
	SIGNAL XSIG825 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X825;
	SIGNAL XSIG826 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X826;
	SIGNAL XSIG827 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X827;
	SIGNAL XSIG828 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X828;
	SIGNAL XSIG829 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X829;
	SIGNAL XSIG830 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X830;
	SIGNAL XSIG831 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X831;
	SIGNAL XSIG832 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X832;
	SIGNAL XSIG833 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X833;
	SIGNAL XSIG834 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X834;
	SIGNAL XSIG835 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X835;
	SIGNAL XSIG836 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X836;
	SIGNAL XSIG837 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X837;
	SIGNAL XSIG838 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X838;
	SIGNAL XSIG839 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X839;
	SIGNAL XSIG840 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X840;
	SIGNAL XSIG841 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X841;
	SIGNAL XSIG842 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X842;
	SIGNAL XSIG843 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X843;
	SIGNAL XSIG844 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X844;
	SIGNAL XSIG845 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X845;
	SIGNAL XSIG846 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X846;
	SIGNAL XSIG847 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X847;
	SIGNAL XSIG848 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X848;
	SIGNAL XSIG849 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X849;
	SIGNAL XSIG850 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X850;
	SIGNAL XSIG851 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X851;
	SIGNAL XSIG852 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X852;
	SIGNAL XSIG853 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X853;
	SIGNAL XSIG854 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X854;
	SIGNAL XSIG855 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X855;
	SIGNAL XSIG856 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X856;
	SIGNAL XSIG857 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X857;
	SIGNAL XSIG858 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X858;
	SIGNAL XSIG859 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X859;
	SIGNAL XSIG860 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X860;
	SIGNAL XSIG861 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X861;
	SIGNAL XSIG862 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X862;
	SIGNAL XSIG863 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X863;
	SIGNAL XSIG864 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X864;
	SIGNAL XSIG865 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X865;
	SIGNAL XSIG866 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X866;
	SIGNAL XSIG867 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X867;
	SIGNAL XSIG868 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X868;
	SIGNAL XSIG869 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X869;
	SIGNAL XSIG870 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X870;
	SIGNAL XSIG871 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X871;
	SIGNAL XSIG872 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X872;
	SIGNAL XSIG873 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X873;
	SIGNAL XSIG874 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X874;
	SIGNAL XSIG875 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X875;
	SIGNAL XSIG876 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X876;
	SIGNAL XSIG877 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X877;
	SIGNAL XSIG878 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X878;
	SIGNAL XSIG879 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X879;
	SIGNAL XSIG880 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X880;
	SIGNAL XSIG881 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X881;
	SIGNAL XSIG882 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X882;
	SIGNAL XSIG883 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X883;
	SIGNAL XSIG884 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X884;
	SIGNAL XSIG885 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X885;
	SIGNAL XSIG886 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X886;
	SIGNAL XSIG887 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X887;
	SIGNAL XSIG888 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X888;
	SIGNAL XSIG889 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X889;
	SIGNAL XSIG890 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X890;
	SIGNAL XSIG891 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X891;
	SIGNAL XSIG892 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X892;
	SIGNAL XSIG893 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X893;
	SIGNAL XSIG894 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X894;
	SIGNAL XSIG895 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X895;
	SIGNAL XSIG896 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X896;
	SIGNAL XSIG897 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X897;
	SIGNAL XSIG898 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X898;
	SIGNAL XSIG899 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X899;
	SIGNAL XSIG900 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X900;
	SIGNAL XSIG901 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X901;
	SIGNAL XSIG902 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X902;
	SIGNAL XSIG903 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X903;
	SIGNAL XSIG904 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X904;
	SIGNAL XSIG905 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X905;
	SIGNAL XSIG906 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X906;
	SIGNAL XSIG907 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X907;
	SIGNAL XSIG908 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X908;
	SIGNAL XSIG909 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X909;
	SIGNAL XSIG910 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X910;
	SIGNAL XSIG911 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X911;
	SIGNAL XSIG912 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X912;
	SIGNAL XSIG913 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X913;
	SIGNAL XSIG914 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X914;
	SIGNAL XSIG915 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X915;
	SIGNAL XSIG916 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X916;
	SIGNAL XSIG917 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X917;
	SIGNAL XSIG918 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X918;
	SIGNAL XSIG919 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X919;
	SIGNAL XSIG920 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X920;
	SIGNAL XSIG921 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X921;
	SIGNAL XSIG922 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X922;
	SIGNAL XSIG923 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X923;
	SIGNAL XSIG924 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X924;
	SIGNAL XSIG925 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X925;
	SIGNAL XSIG926 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X926;
	SIGNAL XSIG927 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X927;
	SIGNAL XSIG928 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X928;
	SIGNAL XSIG929 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X929;
	SIGNAL XSIG930 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X930;
	SIGNAL XSIG931 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X931;
	SIGNAL XSIG932 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X932;
	SIGNAL XSIG933 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X933;
	SIGNAL XSIG934 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X934;
	SIGNAL XSIG935 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X935;
	SIGNAL XSIG936 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X936;
	SIGNAL XSIG937 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X937;
	SIGNAL XSIG938 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X938;
	SIGNAL XSIG939 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X939;
	SIGNAL XSIG940 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X940;
	SIGNAL XSIG941 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X941;
	SIGNAL XSIG942 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X942;
	SIGNAL XSIG943 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X943;
	SIGNAL XSIG944 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X944;
	SIGNAL XSIG945 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X945;
	SIGNAL XSIG946 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X946;
	SIGNAL XSIG947 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X947;
	SIGNAL XSIG948 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X948;
	SIGNAL XSIG949 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X949;
	SIGNAL XSIG950 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X950;
	SIGNAL XSIG951 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X951;
	SIGNAL XSIG952 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X952;
	SIGNAL XSIG953 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X953;
	SIGNAL XSIG954 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X954;
	SIGNAL XSIG955 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X955;
	SIGNAL XSIG956 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X956;
	SIGNAL XSIG957 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X957;
	SIGNAL XSIG958 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X958;
	SIGNAL XSIG959 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X959;
	SIGNAL XSIG960 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X960;
	SIGNAL XSIG961 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X961;
	SIGNAL XSIG962 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X962;
	SIGNAL XSIG963 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X963;
	SIGNAL XSIG964 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X964;
	SIGNAL XSIG965 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X965;
	SIGNAL XSIG966 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X966;
	SIGNAL XSIG967 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X967;
	SIGNAL XSIG968 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X968;
	SIGNAL XSIG969 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X969;
	SIGNAL XSIG970 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X970;
	SIGNAL XSIG971 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X971;
	SIGNAL XSIG972 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X972;
	SIGNAL XSIG973 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X973;
	SIGNAL XSIG974 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X974;
	SIGNAL XSIG975 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X975;
	SIGNAL XSIG976 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X976;
	SIGNAL XSIG977 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X977;
	SIGNAL XSIG978 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X978;
	SIGNAL XSIG979 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X979;
	SIGNAL XSIG980 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X980;
	SIGNAL XSIG981 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X981;
	SIGNAL XSIG982 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X982;
	SIGNAL XSIG983 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X983;
	SIGNAL XSIG984 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X984;
	SIGNAL XSIG985 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X985;
	SIGNAL XSIG986 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X986;
	SIGNAL XSIG987 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X987;
	SIGNAL XSIG988 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X988;
	SIGNAL XSIG989 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X989;
	SIGNAL XSIG990 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X990;
	SIGNAL XSIG991 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X991;
	SIGNAL XSIG992 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X992;
	SIGNAL XSIG993 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X993;
	SIGNAL XSIG994 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X994;
	SIGNAL XSIG995 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X995;
	SIGNAL XSIG996 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X996;
	SIGNAL XSIG997 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X997;
	SIGNAL XSIG998 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X998;
	SIGNAL XSIG999 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X999;
	SIGNAL XSIG1000 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1000;
	SIGNAL XSIG1001 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1001;
	SIGNAL XSIG1002 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1002;
	SIGNAL XSIG1003 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1003;
	SIGNAL XSIG1004 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1004;
	SIGNAL XSIG1005 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1005;
	SIGNAL XSIG1006 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1006;
	SIGNAL XSIG1007 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1007;
	SIGNAL XSIG1008 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1008;
	SIGNAL XSIG1009 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1009;
	SIGNAL XSIG1010 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1010;
	SIGNAL XSIG1011 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1011;
	SIGNAL XSIG1012 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1012;
	SIGNAL XSIG1013 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1013;
	SIGNAL XSIG1014 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1014;
	SIGNAL XSIG1015 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1015;
	SIGNAL XSIG1016 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1016;
	SIGNAL XSIG1017 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1017;
	SIGNAL XSIG1018 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1018;
	SIGNAL XSIG1019 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1019;
	SIGNAL XSIG1020 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1020;
	SIGNAL XSIG1021 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1021;
	SIGNAL XSIG1022 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1022;
	SIGNAL XSIG1023 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1023;
	SIGNAL XSIG1024 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1024;
	SIGNAL XSIG1025 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1025;
	SIGNAL XSIG1026 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1026;
	SIGNAL XSIG1027 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1027;
	SIGNAL XSIG1028 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1028;
	SIGNAL XSIG1029 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1029;
	SIGNAL XSIG1030 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1030;
	SIGNAL XSIG1031 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1031;
	SIGNAL XSIG1032 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1032;
	SIGNAL XSIG1033 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1033;
	SIGNAL XSIG1034 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1034;
	SIGNAL XSIG1035 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1035;
	SIGNAL XSIG1036 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1036;
	SIGNAL XSIG1037 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1037;
	SIGNAL XSIG1038 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1038;
	SIGNAL XSIG1039 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1039;
	SIGNAL XSIG1040 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1040;
	SIGNAL XSIG1041 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1041;
	SIGNAL XSIG1042 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1042;
	SIGNAL XSIG1043 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1043;
	SIGNAL XSIG1044 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1044;
	SIGNAL XSIG1045 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1045;
	SIGNAL XSIG1046 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1046;
	SIGNAL XSIG1047 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1047;
	SIGNAL XSIG1048 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1048;
	SIGNAL XSIG1049 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1049;
	SIGNAL XSIG1050 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1050;
	SIGNAL XSIG1051 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1051;
	SIGNAL XSIG1052 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1052;
	SIGNAL XSIG1053 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1053;
	SIGNAL XSIG1054 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1054;
	SIGNAL XSIG1055 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1055;
	SIGNAL XSIG1056 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1056;
	SIGNAL XSIG1057 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1057;
	SIGNAL XSIG1058 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1058;
	SIGNAL XSIG1059 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1059;
	SIGNAL XSIG1060 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1060;
	SIGNAL XSIG1061 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1061;
	SIGNAL XSIG1062 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1062;
	SIGNAL XSIG1063 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1063;
	SIGNAL XSIG1064 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1064;
	SIGNAL XSIG1065 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1065;
	SIGNAL XSIG1066 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1066;
	SIGNAL XSIG1067 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1067;
	SIGNAL XSIG1068 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1068;
	SIGNAL XSIG1069 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1069;
	SIGNAL XSIG1070 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1070;
	SIGNAL XSIG1071 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1071;
	SIGNAL XSIG1072 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1072;
	SIGNAL XSIG1073 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1073;
	SIGNAL XSIG1074 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1074;
	SIGNAL XSIG1075 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1075;
	SIGNAL XSIG1076 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1076;
	SIGNAL XSIG1077 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1077;
	SIGNAL XSIG1078 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1078;
	SIGNAL XSIG1079 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1079;
	SIGNAL XSIG1080 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1080;
	SIGNAL XSIG1081 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1081;
	SIGNAL XSIG1082 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1082;
	SIGNAL XSIG1083 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1083;
	SIGNAL XSIG1084 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1084;
	SIGNAL XSIG1085 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1085;
	SIGNAL XSIG1086 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1086;
	SIGNAL XSIG1087 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1087;
	SIGNAL XSIG1088 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1088;
	SIGNAL XSIG1089 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1089;
	SIGNAL XSIG1090 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1090;
	SIGNAL XSIG1091 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1091;
	SIGNAL XSIG1092 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1092;
	SIGNAL XSIG1093 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1093;
	SIGNAL XSIG1094 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1094;
	SIGNAL XSIG1095 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1095;
	SIGNAL XSIG1096 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1096;
	SIGNAL XSIG1097 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1097;
	SIGNAL XSIG1098 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1098;
	SIGNAL XSIG1099 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1099;
	SIGNAL XSIG1100 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1100;
	SIGNAL XSIG1101 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1101;
	SIGNAL XSIG1102 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1102;
	SIGNAL XSIG1103 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1103;
	SIGNAL XSIG1104 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1104;
	SIGNAL XSIG1105 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1105;
	SIGNAL XSIG1106 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1106;
	SIGNAL XSIG1107 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1107;
	SIGNAL XSIG1108 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1108;
	SIGNAL XSIG1109 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1109;
	SIGNAL XSIG1110 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1110;
	SIGNAL XSIG1111 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1111;
	SIGNAL XSIG1112 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1112;
	SIGNAL XSIG1113 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1113;
	SIGNAL XSIG1114 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1114;
	SIGNAL XSIG1115 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1115;
	SIGNAL XSIG1116 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1116;
	SIGNAL XSIG1117 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1117;
	SIGNAL XSIG1118 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1118;
	SIGNAL XSIG1119 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1119;
	SIGNAL XSIG1120 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1120;
	SIGNAL XSIG1121 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1121;
	SIGNAL XSIG1122 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1122;
	SIGNAL XSIG1123 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1123;
	SIGNAL XSIG1124 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1124;
	SIGNAL XSIG1125 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1125;
	SIGNAL XSIG1126 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1126;
	SIGNAL XSIG1127 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1127;
	SIGNAL XSIG1128 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1128;
	SIGNAL XSIG1129 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1129;
	SIGNAL XSIG1130 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1130;
	SIGNAL XSIG1131 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1131;
	SIGNAL XSIG1132 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1132;
	SIGNAL XSIG1133 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1133;
	SIGNAL XSIG1134 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1134;
	SIGNAL XSIG1135 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1135;
	SIGNAL XSIG1136 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1136;
	SIGNAL XSIG1137 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1137;
	SIGNAL XSIG1138 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1138;
	SIGNAL XSIG1139 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1139;
	SIGNAL XSIG1140 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1140;
	SIGNAL XSIG1141 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1141;
	SIGNAL XSIG1142 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1142;
	SIGNAL XSIG1143 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1143;
	SIGNAL XSIG1144 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1144;
	SIGNAL XSIG1145 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1145;
	SIGNAL XSIG1146 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1146;
	SIGNAL XSIG1147 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1147;
	SIGNAL XSIG1148 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1148;
	SIGNAL XSIG1149 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1149;
	SIGNAL XSIG1150 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1150;
	SIGNAL XSIG1151 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1151;
	SIGNAL XSIG1152 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1152;
	SIGNAL XSIG1153 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1153;
	SIGNAL XSIG1154 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1154;
	SIGNAL XSIG1155 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1155;
	SIGNAL XSIG1156 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1156;
	SIGNAL XSIG1157 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1157;
	SIGNAL XSIG1158 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1158;
	SIGNAL XSIG1159 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1159;
	SIGNAL XSIG1160 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1160;
	SIGNAL XSIG1161 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1161;
	SIGNAL XSIG1162 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1162;
	SIGNAL XSIG1163 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1163;
	SIGNAL XSIG1164 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1164;
	SIGNAL XSIG1165 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1165;
	SIGNAL XSIG1166 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1166;
	SIGNAL XSIG1167 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1167;
	SIGNAL XSIG1168 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1168;
	SIGNAL XSIG1169 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1169;
	SIGNAL XSIG1170 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1170;
	SIGNAL XSIG1171 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1171;
	SIGNAL XSIG1172 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1172;
	SIGNAL XSIG1173 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1173;
	SIGNAL XSIG1174 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1174;
	SIGNAL XSIG1175 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1175;
	SIGNAL XSIG1176 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1176;
	SIGNAL XSIG1177 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1177;
	SIGNAL XSIG1178 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1178;
	SIGNAL XSIG1179 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1179;
	SIGNAL XSIG1180 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1180;
	SIGNAL XSIG1181 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1181;
	SIGNAL XSIG1182 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1182;
	SIGNAL XSIG1183 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1183;
	SIGNAL XSIG1184 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1184;
	SIGNAL XSIG1185 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1185;
	SIGNAL XSIG1186 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1186;
	SIGNAL XSIG1187 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1187;
	SIGNAL XSIG1188 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1188;
	SIGNAL XSIG1189 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1189;
	SIGNAL XSIG1190 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1190;
	SIGNAL XSIG1191 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1191;
	SIGNAL XSIG1192 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1192;
	SIGNAL XSIG1193 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1193;
	SIGNAL XSIG1194 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1194;
	SIGNAL XSIG1195 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1195;
	SIGNAL XSIG1196 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1196;
	SIGNAL XSIG1197 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1197;
	SIGNAL XSIG1198 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1198;
	SIGNAL XSIG1199 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1199;
	SIGNAL XSIG1200 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1200;
	SIGNAL XSIG1201 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1201;
	SIGNAL XSIG1202 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1202;
	SIGNAL XSIG1203 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1203;
	SIGNAL XSIG1204 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1204;
	SIGNAL XSIG1205 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1205;
	SIGNAL XSIG1206 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1206;
	SIGNAL XSIG1207 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1207;
	SIGNAL XSIG1208 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1208;
	SIGNAL XSIG1209 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1209;
	SIGNAL XSIG1210 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1210;
	SIGNAL XSIG1211 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1211;
	SIGNAL XSIG1212 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1212;
	SIGNAL XSIG1213 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1213;
	SIGNAL XSIG1214 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1214;
	SIGNAL XSIG1215 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1215;
	SIGNAL XSIG1216 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1216;
	SIGNAL XSIG1217 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1217;
	SIGNAL XSIG1218 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1218;
	SIGNAL XSIG1219 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1219;
	SIGNAL XSIG1220 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1220;
	SIGNAL XSIG1221 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1221;
	SIGNAL XSIG1222 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1222;
	SIGNAL XSIG1223 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1223;
	SIGNAL XSIG1224 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1224;
	SIGNAL XSIG1225 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1225;
	SIGNAL XSIG1226 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1226;
	SIGNAL XSIG1227 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1227;
	SIGNAL XSIG1228 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1228;
	SIGNAL XSIG1229 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1229;
	SIGNAL XSIG1230 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1230;
	SIGNAL XSIG1231 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1231;
	SIGNAL XSIG1232 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1232;
	SIGNAL XSIG1233 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1233;
	SIGNAL XSIG1234 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1234;
	SIGNAL XSIG1235 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1235;
	SIGNAL XSIG1236 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1236;
	SIGNAL XSIG1237 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1237;
	SIGNAL XSIG1238 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1238;
	SIGNAL XSIG1239 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1239;
	SIGNAL XSIG1240 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1240;
	SIGNAL XSIG1241 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1241;
	SIGNAL XSIG1242 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1242;
	SIGNAL XSIG1243 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1243;
	SIGNAL XSIG1244 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1244;
	SIGNAL XSIG1245 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1245;
	SIGNAL XSIG1246 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1246;
	SIGNAL XSIG1247 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1247;
	SIGNAL XSIG1248 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1248;
	SIGNAL XSIG1249 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1249;
	SIGNAL XSIG1250 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1250;
	SIGNAL XSIG1251 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1251;
	SIGNAL XSIG1252 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1252;
	SIGNAL XSIG1253 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1253;
	SIGNAL XSIG1254 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1254;
	SIGNAL XSIG1255 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1255;
	SIGNAL XSIG1256 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1256;
	SIGNAL XSIG1257 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1257;
	SIGNAL XSIG1258 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1258;
	SIGNAL XSIG1259 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1259;
	SIGNAL XSIG1260 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1260;
	SIGNAL XSIG1261 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1261;
	SIGNAL XSIG1262 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1262;
	SIGNAL XSIG1263 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1263;
	SIGNAL XSIG1264 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1264;
	SIGNAL XSIG1265 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1265;
	SIGNAL XSIG1266 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1266;
	SIGNAL XSIG1267 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1267;
	SIGNAL XSIG1268 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1268;
	SIGNAL XSIG1269 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1269;
	SIGNAL XSIG1270 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1270;
	SIGNAL XSIG1271 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1271;
	SIGNAL XSIG1272 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1272;
	SIGNAL XSIG1273 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1273;
	SIGNAL XSIG1274 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1274;
	SIGNAL XSIG1275 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1275;
	SIGNAL XSIG1276 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1276;
	SIGNAL XSIG1277 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1277;
	SIGNAL XSIG1278 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1278;
	SIGNAL XSIG1279 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1279;
	SIGNAL XSIG1280 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1280;
	SIGNAL XSIG1281 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1281;
	SIGNAL XSIG1282 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1282;
	SIGNAL XSIG1283 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1283;
	SIGNAL XSIG1284 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1284;
	SIGNAL XSIG1285 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1285;
	SIGNAL XSIG1286 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1286;
	SIGNAL XSIG1287 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1287;
	SIGNAL XSIG1288 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1288;
	SIGNAL XSIG1289 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1289;
	SIGNAL XSIG1290 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1290;
	SIGNAL XSIG1291 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1291;
	SIGNAL XSIG1292 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1292;
	SIGNAL XSIG1293 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1293;
	SIGNAL XSIG1294 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1294;
	SIGNAL XSIG1295 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1295;
	SIGNAL XSIG1296 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1296;
	SIGNAL XSIG1297 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1297;
	SIGNAL XSIG1298 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1298;
	SIGNAL XSIG1299 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1299;
	SIGNAL XSIG1300 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1300;
	SIGNAL XSIG1301 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1301;
	SIGNAL XSIG1302 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1302;
	SIGNAL XSIG1303 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1303;
	SIGNAL XSIG1304 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1304;
	SIGNAL XSIG1305 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1305;
	SIGNAL XSIG1306 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1306;
	SIGNAL XSIG1307 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1307;
	SIGNAL XSIG1308 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1308;
	SIGNAL XSIG1309 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1309;
	SIGNAL XSIG1310 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1310;
	SIGNAL XSIG1311 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1311;
	SIGNAL XSIG1312 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1312;
	SIGNAL XSIG1313 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1313;
	SIGNAL XSIG1314 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1314;
	SIGNAL XSIG1315 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1315;
	SIGNAL XSIG1316 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1316;
	SIGNAL XSIG1317 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1317;
	SIGNAL XSIG1318 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1318;
	SIGNAL XSIG1319 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1319;
	SIGNAL XSIG1320 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1320;
	SIGNAL XSIG1321 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1321;
	SIGNAL XSIG1322 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1322;
	SIGNAL XSIG1323 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1323;
	SIGNAL XSIG1324 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1324;
	SIGNAL XSIG1325 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1325;
	SIGNAL XSIG1326 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1326;
	SIGNAL XSIG1327 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1327;
	SIGNAL XSIG1328 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1328;
	SIGNAL XSIG1329 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1329;
	SIGNAL XSIG1330 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1330;
	SIGNAL XSIG1331 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1331;
	SIGNAL XSIG1332 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1332;
	SIGNAL XSIG1333 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1333;
	SIGNAL XSIG1334 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1334;
	SIGNAL XSIG1335 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1335;
	SIGNAL XSIG1336 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1336;
	SIGNAL XSIG1337 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1337;
	SIGNAL XSIG1338 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1338;
	SIGNAL XSIG1339 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1339;
	SIGNAL XSIG1340 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1340;
	SIGNAL XSIG1341 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1341;
	SIGNAL XSIG1342 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1342;
	SIGNAL XSIG1343 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1343;
	SIGNAL XSIG1344 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1344;
	SIGNAL XSIG1345 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1345;
	SIGNAL XSIG1346 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1346;
	SIGNAL XSIG1347 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1347;
	SIGNAL XSIG1348 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1348;
	SIGNAL XSIG1349 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1349;
	SIGNAL XSIG1350 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1350;
	SIGNAL XSIG1351 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1351;
	SIGNAL XSIG1352 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1352;
	SIGNAL XSIG1353 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1353;
	SIGNAL XSIG1354 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1354;
	SIGNAL XSIG1355 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1355;
	SIGNAL XSIG1356 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1356;
	SIGNAL XSIG1357 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1357;
	SIGNAL XSIG1358 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1358;
	SIGNAL XSIG1359 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1359;
	SIGNAL XSIG1360 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1360;
	SIGNAL XSIG1361 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1361;
	SIGNAL XSIG1362 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1362;
	SIGNAL XSIG1363 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1363;
	SIGNAL XSIG1364 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1364;
	SIGNAL XSIG1365 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1365;
	SIGNAL XSIG1366 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1366;
	SIGNAL XSIG1367 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1367;
	SIGNAL XSIG1368 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1368;
	SIGNAL XSIG1369 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1369;
	SIGNAL XSIG1370 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1370;
	SIGNAL XSIG1371 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1371;
	SIGNAL XSIG1372 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1372;
	SIGNAL XSIG1373 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1373;
	SIGNAL XSIG1374 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1374;
	SIGNAL XSIG1375 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1375;
	SIGNAL XSIG1376 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1376;
	SIGNAL XSIG1377 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1377;
	SIGNAL XSIG1378 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1378;
	SIGNAL XSIG1379 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1379;
	SIGNAL XSIG1380 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1380;
	SIGNAL XSIG1381 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1381;
	SIGNAL XSIG1382 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1382;
	SIGNAL XSIG1383 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1383;
	SIGNAL XSIG1384 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1384;
	SIGNAL XSIG1385 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1385;
	SIGNAL XSIG1386 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1386;
	SIGNAL XSIG1387 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1387;
	SIGNAL XSIG1388 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1388;
	SIGNAL XSIG1389 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1389;
	SIGNAL XSIG1390 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1390;
	SIGNAL XSIG1391 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1391;
	SIGNAL XSIG1392 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1392;
	SIGNAL XSIG1393 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1393;
	SIGNAL XSIG1394 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1394;
	SIGNAL XSIG1395 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1395;
	SIGNAL XSIG1396 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1396;
	SIGNAL XSIG1397 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1397;
	SIGNAL XSIG1398 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1398;
	SIGNAL XSIG1399 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1399;
	SIGNAL XSIG1400 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1400;
	SIGNAL XSIG1401 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1401;
	SIGNAL XSIG1402 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1402;
	SIGNAL XSIG1403 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1403;
	SIGNAL XSIG1404 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1404;
	SIGNAL XSIG1405 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1405;
	SIGNAL XSIG1406 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1406;
	SIGNAL XSIG1407 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1407;
	SIGNAL XSIG1408 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1408;
	SIGNAL XSIG1409 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1409;
	SIGNAL XSIG1410 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1410;
	SIGNAL XSIG1411 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1411;
	SIGNAL XSIG1412 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1412;
	SIGNAL XSIG1413 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1413;
	SIGNAL XSIG1414 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1414;
	SIGNAL XSIG1415 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1415;
	SIGNAL XSIG1416 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1416;
	SIGNAL XSIG1417 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1417;
	SIGNAL XSIG1418 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1418;
	SIGNAL XSIG1419 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1419;
	SIGNAL XSIG1420 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1420;
	SIGNAL XSIG1421 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1421;
	SIGNAL XSIG1422 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1422;
	SIGNAL XSIG1423 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1423;
	SIGNAL XSIG1424 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1424;
	SIGNAL XSIG1425 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1425;
	SIGNAL XSIG1426 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1426;
	SIGNAL XSIG1427 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1427;
	SIGNAL XSIG1428 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1428;
	SIGNAL XSIG1429 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1429;
	SIGNAL XSIG1430 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1430;
	SIGNAL XSIG1431 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1431;
	SIGNAL XSIG1432 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1432;
	SIGNAL XSIG1433 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1433;
	SIGNAL XSIG1434 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1434;
	SIGNAL XSIG1435 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1435;
	SIGNAL XSIG1436 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1436;
	SIGNAL XSIG1437 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1437;
	SIGNAL XSIG1438 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1438;
	SIGNAL XSIG1439 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1439;
	SIGNAL XSIG1440 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1440;
	SIGNAL XSIG1441 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1441;
	SIGNAL XSIG1442 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1442;
	SIGNAL XSIG1443 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1443;
	SIGNAL XSIG1444 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1444;
	SIGNAL XSIG1445 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1445;
	SIGNAL XSIG1446 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1446;
	SIGNAL XSIG1447 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1447;
	SIGNAL XSIG1448 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1448;
	SIGNAL XSIG1449 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1449;
	SIGNAL XSIG1450 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1450;
	SIGNAL XSIG1451 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1451;
	SIGNAL XSIG1452 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1452;
	SIGNAL XSIG1453 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1453;
	SIGNAL XSIG1454 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1454;
	SIGNAL XSIG1455 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1455;
	SIGNAL XSIG1456 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1456;
	SIGNAL XSIG1457 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1457;
	SIGNAL XSIG1458 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1458;
	SIGNAL XSIG1459 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1459;
	SIGNAL XSIG1460 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1460;
	SIGNAL XSIG1461 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1461;
	SIGNAL XSIG1462 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1462;
	SIGNAL XSIG1463 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1463;
	SIGNAL XSIG1464 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1464;
	SIGNAL XSIG1465 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1465;
	SIGNAL XSIG1466 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1466;
	SIGNAL XSIG1467 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1467;
	SIGNAL XSIG1468 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1468;
	SIGNAL XSIG1469 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1469;
	SIGNAL XSIG1470 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1470;
	SIGNAL XSIG1471 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1471;
	SIGNAL XSIG1472 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1472;
	SIGNAL XSIG1473 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1473;
	SIGNAL XSIG1474 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1474;
	SIGNAL XSIG1475 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1475;
	SIGNAL XSIG1476 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1476;
	SIGNAL XSIG1477 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1477;
	SIGNAL XSIG1478 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1478;
	SIGNAL XSIG1479 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1479;
	SIGNAL XSIG1480 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1480;
	SIGNAL XSIG1481 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1481;
	SIGNAL XSIG1482 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1482;
	SIGNAL XSIG1483 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1483;
	SIGNAL XSIG1484 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1484;
	SIGNAL XSIG1485 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1485;
	SIGNAL XSIG1486 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1486;
	SIGNAL XSIG1487 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1487;
	SIGNAL XSIG1488 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1488;
	SIGNAL XSIG1489 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1489;
	SIGNAL XSIG1490 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1490;
	SIGNAL XSIG1491 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1491;
	SIGNAL XSIG1492 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1492;
	SIGNAL XSIG1493 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1493;
	SIGNAL XSIG1494 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1494;
	SIGNAL XSIG1495 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1495;
	SIGNAL XSIG1496 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1496;
	SIGNAL XSIG1497 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1497;
	SIGNAL XSIG1498 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1498;
	SIGNAL XSIG1499 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1499;
	SIGNAL XSIG1500 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1500;
	SIGNAL XSIG1501 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1501;
	SIGNAL XSIG1502 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1502;
	SIGNAL XSIG1503 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1503;
	SIGNAL XSIG1504 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1504;
	SIGNAL XSIG1505 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1505;
	SIGNAL XSIG1506 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1506;
	SIGNAL XSIG1507 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1507;
	SIGNAL XSIG1508 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1508;
	SIGNAL XSIG1509 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1509;
	SIGNAL XSIG1510 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1510;
	SIGNAL XSIG1511 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1511;
	SIGNAL XSIG1512 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1512;
	SIGNAL XSIG1513 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1513;
	SIGNAL XSIG1514 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1514;
	SIGNAL XSIG1515 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1515;
	SIGNAL XSIG1516 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1516;
	SIGNAL XSIG1517 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1517;
	SIGNAL XSIG1518 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1518;
	SIGNAL XSIG1519 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1519;
	SIGNAL XSIG1520 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1520;
	SIGNAL XSIG1521 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1521;
	SIGNAL XSIG1522 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1522;
	SIGNAL XSIG1523 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1523;
	SIGNAL XSIG1524 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1524;
	SIGNAL XSIG1525 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1525;
	SIGNAL XSIG1526 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1526;
	SIGNAL XSIG1527 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1527;
	SIGNAL XSIG1528 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1528;
	SIGNAL XSIG1529 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1529;
	SIGNAL XSIG1530 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1530;
	SIGNAL XSIG1531 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1531;
	SIGNAL XSIG1532 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1532;
	SIGNAL XSIG1533 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1533;
	SIGNAL XSIG1534 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1534;
	SIGNAL XSIG1535 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1535;
	SIGNAL XSIG1536 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1536;
	SIGNAL XSIG1537 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1537;
	SIGNAL XSIG1538 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1538;
	SIGNAL XSIG1539 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1539;
	SIGNAL XSIG1540 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1540;
	SIGNAL XSIG1541 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1541;
	SIGNAL XSIG1542 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1542;
	SIGNAL XSIG1543 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1543;
	SIGNAL XSIG1544 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1544;
	SIGNAL XSIG1545 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1545;
	SIGNAL XSIG1546 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1546;
	SIGNAL XSIG1547 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1547;
	SIGNAL XSIG1548 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1548;
	SIGNAL XSIG1549 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1549;
	SIGNAL XSIG1550 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1550;
	SIGNAL XSIG1551 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1551;
	SIGNAL XSIG1552 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1552;
	SIGNAL XSIG1553 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1553;
	SIGNAL XSIG1554 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1554;
	SIGNAL XSIG1555 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1555;
	SIGNAL XSIG1556 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1556;
	SIGNAL XSIG1557 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1557;
	SIGNAL XSIG1558 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1558;
	SIGNAL XSIG1559 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1559;
	SIGNAL XSIG1560 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1560;
	SIGNAL XSIG1561 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1561;
	SIGNAL XSIG1562 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1562;
	SIGNAL XSIG1563 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1563;
	SIGNAL XSIG1564 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1564;
	SIGNAL XSIG1565 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1565;
	SIGNAL XSIG1566 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1566;
	SIGNAL XSIG1567 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1567;
	SIGNAL XSIG1568 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1568;
	SIGNAL XSIG1569 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1569;
	SIGNAL XSIG1570 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1570;
	SIGNAL XSIG1571 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1571;
	SIGNAL XSIG1572 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1572;
	SIGNAL XSIG1573 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1573;
	SIGNAL XSIG1574 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1574;
	SIGNAL XSIG1575 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1575;
	SIGNAL XSIG1576 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1576;
	SIGNAL XSIG1577 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1577;
	SIGNAL XSIG1578 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1578;
	SIGNAL XSIG1579 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1579;
	SIGNAL XSIG1580 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1580;
	SIGNAL XSIG1581 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1581;
	SIGNAL XSIG1582 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1582;
	SIGNAL XSIG1583 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1583;
	SIGNAL XSIG1584 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1584;
	SIGNAL XSIG1585 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1585;
	SIGNAL XSIG1586 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1586;
	SIGNAL XSIG1587 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1587;
	SIGNAL XSIG1588 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1588;
	SIGNAL XSIG1589 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1589;
	SIGNAL XSIG1590 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1590;
	SIGNAL XSIG1591 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1591;
	SIGNAL XSIG1592 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1592;
	SIGNAL XSIG1593 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1593;
	SIGNAL XSIG1594 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1594;
	SIGNAL XSIG1595 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1595;
	SIGNAL XSIG1596 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1596;
	SIGNAL XSIG1597 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1597;
	SIGNAL XSIG1598 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1598;
	SIGNAL XSIG1599 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1599;
	SIGNAL XSIG1600 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1600;
	SIGNAL XSIG1601 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1601;
	SIGNAL XSIG1602 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1602;
	SIGNAL XSIG1603 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1603;
	SIGNAL XSIG1604 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1604;
	SIGNAL XSIG1605 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1605;
	SIGNAL XSIG1606 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1606;
	SIGNAL XSIG1607 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1607;
	SIGNAL XSIG1608 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1608;
	SIGNAL XSIG1609 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1609;
	SIGNAL XSIG1610 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1610;
	SIGNAL XSIG1611 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1611;
	SIGNAL XSIG1612 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1612;
	SIGNAL XSIG1613 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1613;
	SIGNAL XSIG1614 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1614;
	SIGNAL XSIG1615 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1615;
	SIGNAL XSIG1616 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1616;
	SIGNAL XSIG1617 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1617;
	SIGNAL XSIG1618 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1618;
	SIGNAL XSIG1619 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1619;
	SIGNAL XSIG1620 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1620;
	SIGNAL XSIG1621 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1621;
	SIGNAL XSIG1622 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1622;
	SIGNAL XSIG1623 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1623;
	SIGNAL XSIG1624 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1624;
	SIGNAL XSIG1625 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1625;
	SIGNAL XSIG1626 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1626;
	SIGNAL XSIG1627 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1627;
	SIGNAL XSIG1628 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1628;
	SIGNAL XSIG1629 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1629;
	SIGNAL XSIG1630 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1630;
	SIGNAL XSIG1631 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1631;
	SIGNAL XSIG1632 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1632;
	SIGNAL XSIG1633 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1633;
	SIGNAL XSIG1634 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1634;
	SIGNAL XSIG1635 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1635;
	SIGNAL XSIG1636 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1636;
	SIGNAL XSIG1637 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1637;
	SIGNAL XSIG1638 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1638;
	SIGNAL XSIG1639 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1639;
	SIGNAL XSIG1640 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1640;
	SIGNAL XSIG1641 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1641;
	SIGNAL XSIG1642 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1642;
	SIGNAL XSIG1643 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1643;
	SIGNAL XSIG1644 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1644;
	SIGNAL XSIG1645 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1645;
	SIGNAL XSIG1646 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1646;
	SIGNAL XSIG1647 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1647;
	SIGNAL XSIG1648 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1648;
	SIGNAL XSIG1649 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1649;
	SIGNAL XSIG1650 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1650;
	SIGNAL XSIG1651 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1651;
	SIGNAL XSIG1652 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1652;
	SIGNAL XSIG1653 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1653;
	SIGNAL XSIG1654 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1654;
	SIGNAL XSIG1655 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1655;
	SIGNAL XSIG1656 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1656;
	SIGNAL XSIG1657 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1657;
	SIGNAL XSIG1658 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1658;
	SIGNAL XSIG1659 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1659;
	SIGNAL XSIG1660 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1660;
	SIGNAL XSIG1661 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1661;
	SIGNAL XSIG1662 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1662;
	SIGNAL XSIG1663 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1663;
	SIGNAL XSIG1664 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1664;
	SIGNAL XSIG1665 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1665;
	SIGNAL XSIG1666 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1666;
	SIGNAL XSIG1667 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1667;
	SIGNAL XSIG1668 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1668;
	SIGNAL XSIG1669 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1669;
	SIGNAL XSIG1670 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1670;
	SIGNAL XSIG1671 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1671;
	SIGNAL XSIG1672 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1672;
	SIGNAL XSIG1673 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1673;
	SIGNAL XSIG1674 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1674;
	SIGNAL XSIG1675 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1675;
	SIGNAL XSIG1676 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1676;
	SIGNAL XSIG1677 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1677;
	SIGNAL XSIG1678 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1678;
	SIGNAL XSIG1679 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1679;
	SIGNAL XSIG1680 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1680;
	SIGNAL XSIG1681 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1681;
	SIGNAL XSIG1682 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1682;
	SIGNAL XSIG1683 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1683;
	SIGNAL XSIG1684 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1684;
	SIGNAL XSIG1685 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1685;
	SIGNAL XSIG1686 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1686;
	SIGNAL XSIG1687 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1687;
	SIGNAL XSIG1688 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1688;
	SIGNAL XSIG1689 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1689;
	SIGNAL XSIG1690 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1690;
	SIGNAL XSIG1691 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1691;
	SIGNAL XSIG1692 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1692;
	SIGNAL XSIG1693 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1693;
	SIGNAL XSIG1694 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1694;
	SIGNAL XSIG1695 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1695;
	SIGNAL XSIG1696 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1696;
	SIGNAL XSIG1697 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1697;
	SIGNAL XSIG1698 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1698;
	SIGNAL XSIG1699 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1699;
	SIGNAL XSIG1700 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1700;
	SIGNAL XSIG1701 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1701;
	SIGNAL XSIG1702 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1702;
	SIGNAL XSIG1703 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1703;
	SIGNAL XSIG1704 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1704;
	SIGNAL XSIG1705 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1705;
	SIGNAL XSIG1706 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1706;
	SIGNAL XSIG1707 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1707;
	SIGNAL XSIG1708 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1708;
	SIGNAL XSIG1709 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1709;
	SIGNAL XSIG1710 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1710;
	SIGNAL XSIG1711 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1711;
	SIGNAL XSIG1712 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1712;
	SIGNAL XSIG1713 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1713;
	SIGNAL XSIG1714 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1714;
	SIGNAL XSIG1715 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1715;
	SIGNAL XSIG1716 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1716;
	SIGNAL XSIG1717 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1717;
	SIGNAL XSIG1718 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1718;
	SIGNAL XSIG1719 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1719;
	SIGNAL XSIG1720 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1720;
	SIGNAL XSIG1721 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1721;
	SIGNAL XSIG1722 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1722;
	SIGNAL XSIG1723 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1723;
	SIGNAL XSIG1724 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1724;
	SIGNAL XSIG1725 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1725;
	SIGNAL XSIG1726 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1726;
	SIGNAL XSIG1727 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1727;
	SIGNAL XSIG1728 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1728;
	SIGNAL XSIG1729 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1729;
	SIGNAL XSIG1730 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1730;
	SIGNAL XSIG1731 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1731;
	SIGNAL XSIG1732 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1732;
	SIGNAL XSIG1733 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1733;
	SIGNAL XSIG1734 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1734;
	SIGNAL XSIG1735 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1735;
	SIGNAL XSIG1736 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1736;
	SIGNAL XSIG1737 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1737;
	SIGNAL XSIG1738 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1738;
	SIGNAL XSIG1739 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1739;
	SIGNAL XSIG1740 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1740;
	SIGNAL XSIG1741 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1741;
	SIGNAL XSIG1742 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1742;
	SIGNAL XSIG1743 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1743;
	SIGNAL XSIG1744 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1744;
	SIGNAL XSIG1745 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1745;
	SIGNAL XSIG1746 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1746;
	SIGNAL XSIG1747 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1747;
	SIGNAL XSIG1748 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1748;
	SIGNAL XSIG1749 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1749;
	SIGNAL XSIG1750 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1750;
	SIGNAL XSIG1751 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1751;
	SIGNAL XSIG1752 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1752;
	SIGNAL XSIG1753 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1753;
	SIGNAL XSIG1754 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1754;
	SIGNAL XSIG1755 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1755;
	SIGNAL XSIG1756 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1756;
	SIGNAL XSIG1757 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1757;
	SIGNAL XSIG1758 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1758;
	SIGNAL XSIG1759 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1759;
	SIGNAL XSIG1760 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1760;
	SIGNAL XSIG1761 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1761;
	SIGNAL XSIG1762 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1762;
	SIGNAL XSIG1763 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1763;
	SIGNAL XSIG1764 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1764;
	SIGNAL XSIG1765 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1765;
	SIGNAL XSIG1766 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1766;
	SIGNAL XSIG1767 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1767;
	SIGNAL XSIG1768 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1768;
	SIGNAL XSIG1769 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1769;
	SIGNAL XSIG1770 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1770;
	SIGNAL XSIG1771 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1771;
	SIGNAL XSIG1772 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1772;
	SIGNAL XSIG1773 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1773;
	SIGNAL XSIG1774 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1774;
	SIGNAL XSIG1775 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1775;
	SIGNAL XSIG1776 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1776;
	SIGNAL XSIG1777 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1777;
	SIGNAL XSIG1778 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1778;
	SIGNAL XSIG1779 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1779;
	SIGNAL XSIG1780 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1780;
	SIGNAL XSIG1781 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1781;
	SIGNAL XSIG1782 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1782;
	SIGNAL XSIG1783 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1783;
	SIGNAL XSIG1784 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1784;
	SIGNAL XSIG1785 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1785;
	SIGNAL XSIG1786 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1786;
	SIGNAL XSIG1787 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1787;
	SIGNAL XSIG1788 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1788;
	SIGNAL XSIG1789 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1789;
	SIGNAL XSIG1790 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1790;
	SIGNAL XSIG1791 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1791;
	SIGNAL XSIG1792 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1792;
	SIGNAL XSIG1793 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1793;
	SIGNAL XSIG1794 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1794;
	SIGNAL XSIG1795 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1795;
	SIGNAL XSIG1796 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1796;
	SIGNAL XSIG1797 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1797;
	SIGNAL XSIG1798 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1798;
	SIGNAL XSIG1799 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1799;
	SIGNAL XSIG1800 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1800;
	SIGNAL XSIG1801 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1801;
	SIGNAL XSIG1802 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1802;
	SIGNAL XSIG1803 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1803;
	SIGNAL XSIG1804 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1804;
	SIGNAL XSIG1805 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1805;
	SIGNAL XSIG1806 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1806;
	SIGNAL XSIG1807 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1807;
	SIGNAL XSIG1808 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1808;
	SIGNAL XSIG1809 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1809;
	SIGNAL XSIG1810 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1810;
	SIGNAL XSIG1811 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1811;
	SIGNAL XSIG1812 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1812;
	SIGNAL XSIG1813 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1813;
	SIGNAL XSIG1814 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1814;
	SIGNAL XSIG1815 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1815;
	SIGNAL XSIG1816 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1816;
	SIGNAL XSIG1817 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1817;
	SIGNAL XSIG1818 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1818;
	SIGNAL XSIG1819 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1819;
	SIGNAL XSIG1820 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1820;
	SIGNAL XSIG1821 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1821;
	SIGNAL XSIG1822 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1822;
	SIGNAL XSIG1823 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1823;
	SIGNAL XSIG1824 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1824;
	SIGNAL XSIG1825 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1825;
	SIGNAL XSIG1826 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1826;
	SIGNAL XSIG1827 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1827;
	SIGNAL XSIG1828 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1828;
	SIGNAL XSIG1829 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1829;
	SIGNAL XSIG1830 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1830;
	SIGNAL XSIG1831 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1831;
	SIGNAL XSIG1832 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1832;
	SIGNAL XSIG1833 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1833;
	SIGNAL XSIG1834 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1834;
	SIGNAL XSIG1835 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1835;
	SIGNAL XSIG1836 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1836;
	SIGNAL XSIG1837 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1837;
	SIGNAL XSIG1838 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1838;
	SIGNAL XSIG1839 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1839;
	SIGNAL XSIG1840 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1840;
	SIGNAL XSIG1841 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1841;
	SIGNAL XSIG1842 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1842;
	SIGNAL XSIG1843 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1843;
	SIGNAL XSIG1844 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1844;
	SIGNAL XSIG1845 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1845;
	SIGNAL XSIG1846 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1846;
	SIGNAL XSIG1847 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1847;
	SIGNAL XSIG1848 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1848;
	SIGNAL XSIG1849 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1849;
	SIGNAL XSIG1850 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1850;
	SIGNAL XSIG1851 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1851;
	SIGNAL XSIG1852 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1852;
	SIGNAL XSIG1853 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1853;
	SIGNAL XSIG1854 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1854;
	SIGNAL XSIG1855 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1855;
	SIGNAL XSIG1856 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1856;
	SIGNAL XSIG1857 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1857;
	SIGNAL XSIG1858 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1858;
	SIGNAL XSIG1859 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1859;
	SIGNAL XSIG1860 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1860;
	SIGNAL XSIG1861 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1861;
	SIGNAL XSIG1862 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1862;
	SIGNAL XSIG1863 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1863;
	SIGNAL XSIG1864 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1864;
	SIGNAL XSIG1865 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1865;
	SIGNAL XSIG1866 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1866;
	SIGNAL XSIG1867 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1867;
	SIGNAL XSIG1868 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1868;
	SIGNAL XSIG1869 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1869;
	SIGNAL XSIG1870 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1870;
	SIGNAL XSIG1871 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1871;
	SIGNAL XSIG1872 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1872;
	SIGNAL XSIG1873 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1873;
	SIGNAL XSIG1874 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1874;
	SIGNAL XSIG1875 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1875;
	SIGNAL XSIG1876 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1876;
	SIGNAL XSIG1877 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1877;
	SIGNAL XSIG1878 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1878;
	SIGNAL XSIG1879 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1879;
	SIGNAL XSIG1880 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1880;
	SIGNAL XSIG1881 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1881;
	SIGNAL XSIG1882 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1882;
	SIGNAL XSIG1883 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1883;
	SIGNAL XSIG1884 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1884;
	SIGNAL XSIG1885 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1885;
	SIGNAL XSIG1886 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1886;
	SIGNAL XSIG1887 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1887;
	SIGNAL XSIG1888 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1888;
	SIGNAL XSIG1889 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1889;
	SIGNAL XSIG1890 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1890;
	SIGNAL XSIG1891 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1891;
	SIGNAL XSIG1892 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1892;
	SIGNAL XSIG1893 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1893;
	SIGNAL XSIG1894 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1894;
	SIGNAL XSIG1895 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1895;
	SIGNAL XSIG1896 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1896;
	SIGNAL XSIG1897 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1897;
	SIGNAL XSIG1898 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1898;
	SIGNAL XSIG1899 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1899;
	SIGNAL XSIG1900 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1900;
	SIGNAL XSIG1901 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1901;
	SIGNAL XSIG1902 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1902;
	SIGNAL XSIG1903 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1903;
	SIGNAL XSIG1904 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1904;
	SIGNAL XSIG1905 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1905;
	SIGNAL XSIG1906 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1906;
	SIGNAL XSIG1907 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1907;
	SIGNAL XSIG1908 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1908;
	SIGNAL XSIG1909 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1909;
	SIGNAL XSIG1910 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1910;
	SIGNAL XSIG1911 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1911;
	SIGNAL XSIG1912 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1912;
	SIGNAL XSIG1913 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1913;
	SIGNAL XSIG1914 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1914;
	SIGNAL XSIG1915 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1915;
	SIGNAL XSIG1916 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1916;
	SIGNAL XSIG1917 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1917;
	SIGNAL XSIG1918 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1918;
	SIGNAL XSIG1919 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1919;
	SIGNAL XSIG1920 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1920;
	SIGNAL XSIG1921 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1921;
	SIGNAL XSIG1922 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1922;
	SIGNAL XSIG1923 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1923;
	SIGNAL XSIG1924 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1924;
	SIGNAL XSIG1925 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1925;
	SIGNAL XSIG1926 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1926;
	SIGNAL XSIG1927 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1927;
	SIGNAL XSIG1928 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1928;
	SIGNAL XSIG1929 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1929;
	SIGNAL XSIG1930 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1930;
	SIGNAL XSIG1931 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1931;
	SIGNAL XSIG1932 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1932;
	SIGNAL XSIG1933 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1933;
	SIGNAL XSIG1934 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1934;
	SIGNAL XSIG1935 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1935;
	SIGNAL XSIG1936 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1936;
	SIGNAL XSIG1937 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1937;
	SIGNAL XSIG1938 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1938;
	SIGNAL XSIG1939 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1939;
	SIGNAL XSIG1940 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1940;
	SIGNAL XSIG1941 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1941;
	SIGNAL XSIG1942 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1942;
	SIGNAL XSIG1943 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1943;
	SIGNAL XSIG1944 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1944;
	SIGNAL XSIG1945 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1945;
	SIGNAL XSIG1946 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1946;
	SIGNAL XSIG1947 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1947;
	SIGNAL XSIG1948 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1948;
	SIGNAL XSIG1949 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1949;
	SIGNAL XSIG1950 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1950;
	SIGNAL XSIG1951 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1951;
	SIGNAL XSIG1952 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1952;
	SIGNAL XSIG1953 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1953;
	SIGNAL XSIG1954 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1954;
	SIGNAL XSIG1955 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1955;
	SIGNAL XSIG1956 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1956;
	SIGNAL XSIG1957 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1957;
	SIGNAL XSIG1958 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1958;
	SIGNAL XSIG1959 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1959;
	SIGNAL XSIG1960 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1960;
	SIGNAL XSIG1961 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1961;
	SIGNAL XSIG1962 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1962;
	SIGNAL XSIG1963 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1963;
	SIGNAL XSIG1964 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1964;
	SIGNAL XSIG1965 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1965;
	SIGNAL XSIG1966 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1966;
	SIGNAL XSIG1967 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1967;
	SIGNAL XSIG1968 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1968;
	SIGNAL XSIG1969 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1969;
	SIGNAL XSIG1970 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1970;
	SIGNAL XSIG1971 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1971;
	SIGNAL XSIG1972 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1972;
	SIGNAL XSIG1973 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1973;
	SIGNAL XSIG1974 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1974;
	SIGNAL XSIG1975 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1975;
	SIGNAL XSIG1976 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1976;
	SIGNAL XSIG1977 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1977;
	SIGNAL XSIG1978 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1978;
	SIGNAL XSIG1979 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1979;
	SIGNAL XSIG1980 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1980;
	SIGNAL XSIG1981 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1981;
	SIGNAL XSIG1982 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1982;
	SIGNAL XSIG1983 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1983;
	SIGNAL XSIG1984 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1984;
	SIGNAL XSIG1985 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1985;
	SIGNAL XSIG1986 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1986;
	SIGNAL XSIG1987 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1987;
	SIGNAL XSIG1988 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1988;
	SIGNAL XSIG1989 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1989;
	SIGNAL XSIG1990 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1990;
	SIGNAL XSIG1991 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1991;
	SIGNAL XSIG1992 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1992;
	SIGNAL XSIG1993 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1993;
	SIGNAL XSIG1994 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1994;
	SIGNAL XSIG1995 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1995;
	SIGNAL XSIG1996 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1996;
	SIGNAL XSIG1997 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1997;
	SIGNAL XSIG1998 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1998;
	SIGNAL XSIG1999 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X1999;
	SIGNAL XSIG2000 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2000;
	SIGNAL XSIG2001 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2001;
	SIGNAL XSIG2002 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2002;
	SIGNAL XSIG2003 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2003;
	SIGNAL XSIG2004 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2004;
	SIGNAL XSIG2005 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2005;
	SIGNAL XSIG2006 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2006;
	SIGNAL XSIG2007 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2007;
	SIGNAL XSIG2008 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2008;
	SIGNAL XSIG2009 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2009;
	SIGNAL XSIG2010 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2010;
	SIGNAL XSIG2011 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2011;
	SIGNAL XSIG2012 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2012;
	SIGNAL XSIG2013 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2013;
	SIGNAL XSIG2014 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2014;
	SIGNAL XSIG2015 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2015;
	SIGNAL XSIG2016 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2016;
	SIGNAL XSIG2017 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2017;
	SIGNAL XSIG2018 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2018;
	SIGNAL XSIG2019 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2019;
	SIGNAL XSIG2020 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2020;
	SIGNAL XSIG2021 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2021;
	SIGNAL XSIG2022 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2022;
	SIGNAL XSIG2023 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2023;
	SIGNAL XSIG2024 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2024;
	SIGNAL XSIG2025 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2025;
	SIGNAL XSIG2026 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2026;
	SIGNAL XSIG2027 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2027;
	SIGNAL XSIG2028 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2028;
	SIGNAL XSIG2029 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2029;
	SIGNAL XSIG2030 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2030;
	SIGNAL XSIG2031 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2031;
	SIGNAL XSIG2032 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2032;
	SIGNAL XSIG2033 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2033;
	SIGNAL XSIG2034 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2034;
	SIGNAL XSIG2035 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2035;
	SIGNAL XSIG2036 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2036;
	SIGNAL XSIG2037 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2037;
	SIGNAL XSIG2038 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2038;
	SIGNAL XSIG2039 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2039;
	SIGNAL XSIG2040 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2040;
	SIGNAL XSIG2041 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2041;
	SIGNAL XSIG2042 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2042;
	SIGNAL XSIG2043 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2043;
	SIGNAL XSIG2044 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2044;
	SIGNAL XSIG2045 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2045;
	SIGNAL XSIG2046 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2046;
	SIGNAL XSIG2047 : STD_LOGIC_VECTOR(9 DOWNTO 0) := X2047;
	
	VARIABLE reading_input : STD_LOGIC := '0';

	--SIGNAL reieving_cows : STD_LOGIC := '0';	-- clocking through 2048 samples flag
	BEGIN

	PROCESS(clk,samples_ready)
		BEGIN
			IF rising_edge(samples_ready) THEN
				reading_input := '1';
			END IF;
			IF rising_edge(FFT_finished) THEN
				reading_input := '0';
			END IF;
			
			IF (reading_input = '1') THEN	-- shift the 2048 samples into the FFT
			--recieving_cows
			IF rising_edge(clk) THEN
					CASE i IS		
					WHEN 0 =>
						shift_out0 <= XSIG0;
						shift_out1 <= XSIG1;
						shift_out2 <= XSIG2;
						shift_out3 <= XSIG3;
						shift_out4 <= XSIG4;
						shift_out5 <= XSIG5;
						shift_out6 <= XSIG6;
						shift_out7 <= XSIG7;
						shift_out8 <= XSIG8;
						shift_out9 <= XSIG9;
						shift_out10 <= XSIG10;
						shift_out11 <= XSIG11;
						shift_out12 <= XSIG12;
						shift_out13 <= XSIG13;
						shift_out14 <= XSIG14;
						shift_out15 <= XSIG15;
						i <= i + 1;
					WHEN 1 =>
						shift_out0 <= XSIG16;
						shift_out1 <= XSIG17;
						shift_out2 <= XSIG18;
						shift_out3 <= XSIG19;
						shift_out4 <= XSIG20;
						shift_out5 <= XSIG21;
						shift_out6 <= XSIG22;
						shift_out7 <= XSIG23;
						shift_out8 <= XSIG24;
						shift_out9 <= XSIG25;
						shift_out10 <= XSIG26;
						shift_out11 <= XSIG27;
						shift_out12 <= XSIG28;
						shift_out13 <= XSIG29;
						shift_out14 <= XSIG30;
						shift_out15 <= XSIG31;
						i <= i + 1;
					WHEN 2 =>
						shift_out0 <= XSIG32;
						shift_out1 <= XSIG33;
						shift_out2 <= XSIG34;
						shift_out3 <= XSIG35;
						shift_out4 <= XSIG36;
						shift_out5 <= XSIG37;
						shift_out6 <= XSIG38;
						shift_out7 <= XSIG39;
						shift_out8 <= XSIG40;
						shift_out9 <= XSIG41;
						shift_out10 <= XSIG42;
						shift_out11 <= XSIG43;
						shift_out12 <= XSIG44;
						shift_out13 <= XSIG45;
						shift_out14 <= XSIG46;
						shift_out15 <= XSIG47;
						i <= i + 1;
					WHEN 3 =>
						shift_out0 <= XSIG48;
						shift_out1 <= XSIG49;
						shift_out2 <= XSIG50;
						shift_out3 <= XSIG51;
						shift_out4 <= XSIG52;
						shift_out5 <= XSIG53;
						shift_out6 <= XSIG54;
						shift_out7 <= XSIG55;
						shift_out8 <= XSIG56;
						shift_out9 <= XSIG57;
						shift_out10 <= XSIG58;
						shift_out11 <= XSIG59;
						shift_out12 <= XSIG60;
						shift_out13 <= XSIG61;
						shift_out14 <= XSIG62;
						shift_out15 <= XSIG63;
						i <= i + 1;
					WHEN 4 =>
						shift_out0 <= XSIG64;
						shift_out1 <= XSIG65;
						shift_out2 <= XSIG66;
						shift_out3 <= XSIG67;
						shift_out4 <= XSIG68;
						shift_out5 <= XSIG69;
						shift_out6 <= XSIG70;
						shift_out7 <= XSIG71;
						shift_out8 <= XSIG72;
						shift_out9 <= XSIG73;
						shift_out10 <= XSIG74;
						shift_out11 <= XSIG75;
						shift_out12 <= XSIG76;
						shift_out13 <= XSIG77;
						shift_out14 <= XSIG78;
						shift_out15 <= XSIG79;
						i <= i + 1;
					WHEN 5 =>
						shift_out0 <= XSIG80;
						shift_out1 <= XSIG81;
						shift_out2 <= XSIG82;
						shift_out3 <= XSIG83;
						shift_out4 <= XSIG84;
						shift_out5 <= XSIG85;
						shift_out6 <= XSIG86;
						shift_out7 <= XSIG87;
						shift_out8 <= XSIG88;
						shift_out9 <= XSIG89;
						shift_out10 <= XSIG90;
						shift_out11 <= XSIG91;
						shift_out12 <= XSIG92;
						shift_out13 <= XSIG93;
						shift_out14 <= XSIG94;
						shift_out15 <= XSIG95;
						i <= i + 1;
					WHEN 6 =>
						shift_out0 <= XSIG96;
						shift_out1 <= XSIG97;
						shift_out2 <= XSIG98;
						shift_out3 <= XSIG99;
						shift_out4 <= XSIG100;
						shift_out5 <= XSIG101;
						shift_out6 <= XSIG102;
						shift_out7 <= XSIG103;
						shift_out8 <= XSIG104;
						shift_out9 <= XSIG105;
						shift_out10 <= XSIG106;
						shift_out11 <= XSIG107;
						shift_out12 <= XSIG108;
						shift_out13 <= XSIG109;
						shift_out14 <= XSIG110;
						shift_out15 <= XSIG111;
						i <= i + 1;
					WHEN 7 =>
						shift_out0 <= XSIG112;
						shift_out1 <= XSIG113;
						shift_out2 <= XSIG114;
						shift_out3 <= XSIG115;
						shift_out4 <= XSIG116;
						shift_out5 <= XSIG117;
						shift_out6 <= XSIG118;
						shift_out7 <= XSIG119;
						shift_out8 <= XSIG120;
						shift_out9 <= XSIG121;
						shift_out10 <= XSIG122;
						shift_out11 <= XSIG123;
						shift_out12 <= XSIG124;
						shift_out13 <= XSIG125;
						shift_out14 <= XSIG126;
						shift_out15 <= XSIG127;
						i <= i + 1;
					WHEN 8 =>
						shift_out0 <= XSIG128;
						shift_out1 <= XSIG129;
						shift_out2 <= XSIG130;
						shift_out3 <= XSIG131;
						shift_out4 <= XSIG132;
						shift_out5 <= XSIG133;
						shift_out6 <= XSIG134;
						shift_out7 <= XSIG135;
						shift_out8 <= XSIG136;
						shift_out9 <= XSIG137;
						shift_out10 <= XSIG138;
						shift_out11 <= XSIG139;
						shift_out12 <= XSIG140;
						shift_out13 <= XSIG141;
						shift_out14 <= XSIG142;
						shift_out15 <= XSIG143;
						i <= i + 1;
					WHEN 9 =>
						shift_out0 <= XSIG144;
						shift_out1 <= XSIG145;
						shift_out2 <= XSIG146;
						shift_out3 <= XSIG147;
						shift_out4 <= XSIG148;
						shift_out5 <= XSIG149;
						shift_out6 <= XSIG150;
						shift_out7 <= XSIG151;
						shift_out8 <= XSIG152;
						shift_out9 <= XSIG153;
						shift_out10 <= XSIG154;
						shift_out11 <= XSIG155;
						shift_out12 <= XSIG156;
						shift_out13 <= XSIG157;
						shift_out14 <= XSIG158;
						shift_out15 <= XSIG159;
						i <= i + 1;
					WHEN 10 =>
						shift_out0 <= XSIG160;
						shift_out1 <= XSIG161;
						shift_out2 <= XSIG162;
						shift_out3 <= XSIG163;
						shift_out4 <= XSIG164;
						shift_out5 <= XSIG165;
						shift_out6 <= XSIG166;
						shift_out7 <= XSIG167;
						shift_out8 <= XSIG168;
						shift_out9 <= XSIG169;
						shift_out10 <= XSIG170;
						shift_out11 <= XSIG171;
						shift_out12 <= XSIG172;
						shift_out13 <= XSIG173;
						shift_out14 <= XSIG174;
						shift_out15 <= XSIG175;
						i <= i + 1;
					WHEN 11 =>
						shift_out0 <= XSIG176;
						shift_out1 <= XSIG177;
						shift_out2 <= XSIG178;
						shift_out3 <= XSIG179;
						shift_out4 <= XSIG180;
						shift_out5 <= XSIG181;
						shift_out6 <= XSIG182;
						shift_out7 <= XSIG183;
						shift_out8 <= XSIG184;
						shift_out9 <= XSIG185;
						shift_out10 <= XSIG186;
						shift_out11 <= XSIG187;
						shift_out12 <= XSIG188;
						shift_out13 <= XSIG189;
						shift_out14 <= XSIG190;
						shift_out15 <= XSIG191;
						i <= i + 1;
					WHEN 12 =>
						shift_out0 <= XSIG192;
						shift_out1 <= XSIG193;
						shift_out2 <= XSIG194;
						shift_out3 <= XSIG195;
						shift_out4 <= XSIG196;
						shift_out5 <= XSIG197;
						shift_out6 <= XSIG198;
						shift_out7 <= XSIG199;
						shift_out8 <= XSIG200;
						shift_out9 <= XSIG201;
						shift_out10 <= XSIG202;
						shift_out11 <= XSIG203;
						shift_out12 <= XSIG204;
						shift_out13 <= XSIG205;
						shift_out14 <= XSIG206;
						shift_out15 <= XSIG207;
						i <= i + 1;
					WHEN 13 =>
						shift_out0 <= XSIG208;
						shift_out1 <= XSIG209;
						shift_out2 <= XSIG210;
						shift_out3 <= XSIG211;
						shift_out4 <= XSIG212;
						shift_out5 <= XSIG213;
						shift_out6 <= XSIG214;
						shift_out7 <= XSIG215;
						shift_out8 <= XSIG216;
						shift_out9 <= XSIG217;
						shift_out10 <= XSIG218;
						shift_out11 <= XSIG219;
						shift_out12 <= XSIG220;
						shift_out13 <= XSIG221;
						shift_out14 <= XSIG222;
						shift_out15 <= XSIG223;
						i <= i + 1;
					WHEN 14 =>
						shift_out0 <= XSIG224;
						shift_out1 <= XSIG225;
						shift_out2 <= XSIG226;
						shift_out3 <= XSIG227;
						shift_out4 <= XSIG228;
						shift_out5 <= XSIG229;
						shift_out6 <= XSIG230;
						shift_out7 <= XSIG231;
						shift_out8 <= XSIG232;
						shift_out9 <= XSIG233;
						shift_out10 <= XSIG234;
						shift_out11 <= XSIG235;
						shift_out12 <= XSIG236;
						shift_out13 <= XSIG237;
						shift_out14 <= XSIG238;
						shift_out15 <= XSIG239;
						i <= i + 1;
					WHEN 15 =>
						shift_out0 <= XSIG240;
						shift_out1 <= XSIG241;
						shift_out2 <= XSIG242;
						shift_out3 <= XSIG243;
						shift_out4 <= XSIG244;
						shift_out5 <= XSIG245;
						shift_out6 <= XSIG246;
						shift_out7 <= XSIG247;
						shift_out8 <= XSIG248;
						shift_out9 <= XSIG249;
						shift_out10 <= XSIG250;
						shift_out11 <= XSIG251;
						shift_out12 <= XSIG252;
						shift_out13 <= XSIG253;
						shift_out14 <= XSIG254;
						shift_out15 <= XSIG255;
						i <= i + 1;
					WHEN 16 =>
						shift_out0 <= XSIG256;
						shift_out1 <= XSIG257;
						shift_out2 <= XSIG258;
						shift_out3 <= XSIG259;
						shift_out4 <= XSIG260;
						shift_out5 <= XSIG261;
						shift_out6 <= XSIG262;
						shift_out7 <= XSIG263;
						shift_out8 <= XSIG264;
						shift_out9 <= XSIG265;
						shift_out10 <= XSIG266;
						shift_out11 <= XSIG267;
						shift_out12 <= XSIG268;
						shift_out13 <= XSIG269;
						shift_out14 <= XSIG270;
						shift_out15 <= XSIG271;
						i <= i + 1;
					WHEN 17 =>
						shift_out0 <= XSIG272;
						shift_out1 <= XSIG273;
						shift_out2 <= XSIG274;
						shift_out3 <= XSIG275;
						shift_out4 <= XSIG276;
						shift_out5 <= XSIG277;
						shift_out6 <= XSIG278;
						shift_out7 <= XSIG279;
						shift_out8 <= XSIG280;
						shift_out9 <= XSIG281;
						shift_out10 <= XSIG282;
						shift_out11 <= XSIG283;
						shift_out12 <= XSIG284;
						shift_out13 <= XSIG285;
						shift_out14 <= XSIG286;
						shift_out15 <= XSIG287;
						i <= i + 1;
					WHEN 18 =>
						shift_out0 <= XSIG288;
						shift_out1 <= XSIG289;
						shift_out2 <= XSIG290;
						shift_out3 <= XSIG291;
						shift_out4 <= XSIG292;
						shift_out5 <= XSIG293;
						shift_out6 <= XSIG294;
						shift_out7 <= XSIG295;
						shift_out8 <= XSIG296;
						shift_out9 <= XSIG297;
						shift_out10 <= XSIG298;
						shift_out11 <= XSIG299;
						shift_out12 <= XSIG300;
						shift_out13 <= XSIG301;
						shift_out14 <= XSIG302;
						shift_out15 <= XSIG303;
						i <= i + 1;
					WHEN 19 =>
						shift_out0 <= XSIG304;
						shift_out1 <= XSIG305;
						shift_out2 <= XSIG306;
						shift_out3 <= XSIG307;
						shift_out4 <= XSIG308;
						shift_out5 <= XSIG309;
						shift_out6 <= XSIG310;
						shift_out7 <= XSIG311;
						shift_out8 <= XSIG312;
						shift_out9 <= XSIG313;
						shift_out10 <= XSIG314;
						shift_out11 <= XSIG315;
						shift_out12 <= XSIG316;
						shift_out13 <= XSIG317;
						shift_out14 <= XSIG318;
						shift_out15 <= XSIG319;
						i <= i + 1;
					WHEN 20 =>
						shift_out0 <= XSIG320;
						shift_out1 <= XSIG321;
						shift_out2 <= XSIG322;
						shift_out3 <= XSIG323;
						shift_out4 <= XSIG324;
						shift_out5 <= XSIG325;
						shift_out6 <= XSIG326;
						shift_out7 <= XSIG327;
						shift_out8 <= XSIG328;
						shift_out9 <= XSIG329;
						shift_out10 <= XSIG330;
						shift_out11 <= XSIG331;
						shift_out12 <= XSIG332;
						shift_out13 <= XSIG333;
						shift_out14 <= XSIG334;
						shift_out15 <= XSIG335;
						i <= i + 1;
					WHEN 21 =>
						shift_out0 <= XSIG336;
						shift_out1 <= XSIG337;
						shift_out2 <= XSIG338;
						shift_out3 <= XSIG339;
						shift_out4 <= XSIG340;
						shift_out5 <= XSIG341;
						shift_out6 <= XSIG342;
						shift_out7 <= XSIG343;
						shift_out8 <= XSIG344;
						shift_out9 <= XSIG345;
						shift_out10 <= XSIG346;
						shift_out11 <= XSIG347;
						shift_out12 <= XSIG348;
						shift_out13 <= XSIG349;
						shift_out14 <= XSIG350;
						shift_out15 <= XSIG351;
						i <= i + 1;
					WHEN 22 =>
						shift_out0 <= XSIG352;
						shift_out1 <= XSIG353;
						shift_out2 <= XSIG354;
						shift_out3 <= XSIG355;
						shift_out4 <= XSIG356;
						shift_out5 <= XSIG357;
						shift_out6 <= XSIG358;
						shift_out7 <= XSIG359;
						shift_out8 <= XSIG360;
						shift_out9 <= XSIG361;
						shift_out10 <= XSIG362;
						shift_out11 <= XSIG363;
						shift_out12 <= XSIG364;
						shift_out13 <= XSIG365;
						shift_out14 <= XSIG366;
						shift_out15 <= XSIG367;
						i <= i + 1;
					WHEN 23 =>
						shift_out0 <= XSIG368;
						shift_out1 <= XSIG369;
						shift_out2 <= XSIG370;
						shift_out3 <= XSIG371;
						shift_out4 <= XSIG372;
						shift_out5 <= XSIG373;
						shift_out6 <= XSIG374;
						shift_out7 <= XSIG375;
						shift_out8 <= XSIG376;
						shift_out9 <= XSIG377;
						shift_out10 <= XSIG378;
						shift_out11 <= XSIG379;
						shift_out12 <= XSIG380;
						shift_out13 <= XSIG381;
						shift_out14 <= XSIG382;
						shift_out15 <= XSIG383;
						i <= i + 1;
					WHEN 24 =>
						shift_out0 <= XSIG384;
						shift_out1 <= XSIG385;
						shift_out2 <= XSIG386;
						shift_out3 <= XSIG387;
						shift_out4 <= XSIG388;
						shift_out5 <= XSIG389;
						shift_out6 <= XSIG390;
						shift_out7 <= XSIG391;
						shift_out8 <= XSIG392;
						shift_out9 <= XSIG393;
						shift_out10 <= XSIG394;
						shift_out11 <= XSIG395;
						shift_out12 <= XSIG396;
						shift_out13 <= XSIG397;
						shift_out14 <= XSIG398;
						shift_out15 <= XSIG399;
						i <= i + 1;
					WHEN 25 =>
						shift_out0 <= XSIG400;
						shift_out1 <= XSIG401;
						shift_out2 <= XSIG402;
						shift_out3 <= XSIG403;
						shift_out4 <= XSIG404;
						shift_out5 <= XSIG405;
						shift_out6 <= XSIG406;
						shift_out7 <= XSIG407;
						shift_out8 <= XSIG408;
						shift_out9 <= XSIG409;
						shift_out10 <= XSIG410;
						shift_out11 <= XSIG411;
						shift_out12 <= XSIG412;
						shift_out13 <= XSIG413;
						shift_out14 <= XSIG414;
						shift_out15 <= XSIG415;
						i <= i + 1;
					WHEN 26 =>
						shift_out0 <= XSIG416;
						shift_out1 <= XSIG417;
						shift_out2 <= XSIG418;
						shift_out3 <= XSIG419;
						shift_out4 <= XSIG420;
						shift_out5 <= XSIG421;
						shift_out6 <= XSIG422;
						shift_out7 <= XSIG423;
						shift_out8 <= XSIG424;
						shift_out9 <= XSIG425;
						shift_out10 <= XSIG426;
						shift_out11 <= XSIG427;
						shift_out12 <= XSIG428;
						shift_out13 <= XSIG429;
						shift_out14 <= XSIG430;
						shift_out15 <= XSIG431;
						i <= i + 1;
					WHEN 27 =>
						shift_out0 <= XSIG432;
						shift_out1 <= XSIG433;
						shift_out2 <= XSIG434;
						shift_out3 <= XSIG435;
						shift_out4 <= XSIG436;
						shift_out5 <= XSIG437;
						shift_out6 <= XSIG438;
						shift_out7 <= XSIG439;
						shift_out8 <= XSIG440;
						shift_out9 <= XSIG441;
						shift_out10 <= XSIG442;
						shift_out11 <= XSIG443;
						shift_out12 <= XSIG444;
						shift_out13 <= XSIG445;
						shift_out14 <= XSIG446;
						shift_out15 <= XSIG447;
						i <= i + 1;
					WHEN 28 =>
						shift_out0 <= XSIG448;
						shift_out1 <= XSIG449;
						shift_out2 <= XSIG450;
						shift_out3 <= XSIG451;
						shift_out4 <= XSIG452;
						shift_out5 <= XSIG453;
						shift_out6 <= XSIG454;
						shift_out7 <= XSIG455;
						shift_out8 <= XSIG456;
						shift_out9 <= XSIG457;
						shift_out10 <= XSIG458;
						shift_out11 <= XSIG459;
						shift_out12 <= XSIG460;
						shift_out13 <= XSIG461;
						shift_out14 <= XSIG462;
						shift_out15 <= XSIG463;
						i <= i + 1;
					WHEN 29 =>
						shift_out0 <= XSIG464;
						shift_out1 <= XSIG465;
						shift_out2 <= XSIG466;
						shift_out3 <= XSIG467;
						shift_out4 <= XSIG468;
						shift_out5 <= XSIG469;
						shift_out6 <= XSIG470;
						shift_out7 <= XSIG471;
						shift_out8 <= XSIG472;
						shift_out9 <= XSIG473;
						shift_out10 <= XSIG474;
						shift_out11 <= XSIG475;
						shift_out12 <= XSIG476;
						shift_out13 <= XSIG477;
						shift_out14 <= XSIG478;
						shift_out15 <= XSIG479;
						i <= i + 1;
					WHEN 30 =>
						shift_out0 <= XSIG480;
						shift_out1 <= XSIG481;
						shift_out2 <= XSIG482;
						shift_out3 <= XSIG483;
						shift_out4 <= XSIG484;
						shift_out5 <= XSIG485;
						shift_out6 <= XSIG486;
						shift_out7 <= XSIG487;
						shift_out8 <= XSIG488;
						shift_out9 <= XSIG489;
						shift_out10 <= XSIG490;
						shift_out11 <= XSIG491;
						shift_out12 <= XSIG492;
						shift_out13 <= XSIG493;
						shift_out14 <= XSIG494;
						shift_out15 <= XSIG495;
						i <= i + 1;
					WHEN 31 =>
						shift_out0 <= XSIG496;
						shift_out1 <= XSIG497;
						shift_out2 <= XSIG498;
						shift_out3 <= XSIG499;
						shift_out4 <= XSIG500;
						shift_out5 <= XSIG501;
						shift_out6 <= XSIG502;
						shift_out7 <= XSIG503;
						shift_out8 <= XSIG504;
						shift_out9 <= XSIG505;
						shift_out10 <= XSIG506;
						shift_out11 <= XSIG507;
						shift_out12 <= XSIG508;
						shift_out13 <= XSIG509;
						shift_out14 <= XSIG510;
						shift_out15 <= XSIG511;
						i <= i + 1;
					WHEN 32 =>
						shift_out0 <= XSIG512;
						shift_out1 <= XSIG513;
						shift_out2 <= XSIG514;
						shift_out3 <= XSIG515;
						shift_out4 <= XSIG516;
						shift_out5 <= XSIG517;
						shift_out6 <= XSIG518;
						shift_out7 <= XSIG519;
						shift_out8 <= XSIG520;
						shift_out9 <= XSIG521;
						shift_out10 <= XSIG522;
						shift_out11 <= XSIG523;
						shift_out12 <= XSIG524;
						shift_out13 <= XSIG525;
						shift_out14 <= XSIG526;
						shift_out15 <= XSIG527;
						i <= i + 1;
					WHEN 33 =>
						shift_out0 <= XSIG528;
						shift_out1 <= XSIG529;
						shift_out2 <= XSIG530;
						shift_out3 <= XSIG531;
						shift_out4 <= XSIG532;
						shift_out5 <= XSIG533;
						shift_out6 <= XSIG534;
						shift_out7 <= XSIG535;
						shift_out8 <= XSIG536;
						shift_out9 <= XSIG537;
						shift_out10 <= XSIG538;
						shift_out11 <= XSIG539;
						shift_out12 <= XSIG540;
						shift_out13 <= XSIG541;
						shift_out14 <= XSIG542;
						shift_out15 <= XSIG543;
						i <= i + 1;
					WHEN 34 =>
						shift_out0 <= XSIG544;
						shift_out1 <= XSIG545;
						shift_out2 <= XSIG546;
						shift_out3 <= XSIG547;
						shift_out4 <= XSIG548;
						shift_out5 <= XSIG549;
						shift_out6 <= XSIG550;
						shift_out7 <= XSIG551;
						shift_out8 <= XSIG552;
						shift_out9 <= XSIG553;
						shift_out10 <= XSIG554;
						shift_out11 <= XSIG555;
						shift_out12 <= XSIG556;
						shift_out13 <= XSIG557;
						shift_out14 <= XSIG558;
						shift_out15 <= XSIG559;
						i <= i + 1;
					WHEN 35 =>
						shift_out0 <= XSIG560;
						shift_out1 <= XSIG561;
						shift_out2 <= XSIG562;
						shift_out3 <= XSIG563;
						shift_out4 <= XSIG564;
						shift_out5 <= XSIG565;
						shift_out6 <= XSIG566;
						shift_out7 <= XSIG567;
						shift_out8 <= XSIG568;
						shift_out9 <= XSIG569;
						shift_out10 <= XSIG570;
						shift_out11 <= XSIG571;
						shift_out12 <= XSIG572;
						shift_out13 <= XSIG573;
						shift_out14 <= XSIG574;
						shift_out15 <= XSIG575;
						i <= i + 1;
					WHEN 36 =>
						shift_out0 <= XSIG576;
						shift_out1 <= XSIG577;
						shift_out2 <= XSIG578;
						shift_out3 <= XSIG579;
						shift_out4 <= XSIG580;
						shift_out5 <= XSIG581;
						shift_out6 <= XSIG582;
						shift_out7 <= XSIG583;
						shift_out8 <= XSIG584;
						shift_out9 <= XSIG585;
						shift_out10 <= XSIG586;
						shift_out11 <= XSIG587;
						shift_out12 <= XSIG588;
						shift_out13 <= XSIG589;
						shift_out14 <= XSIG590;
						shift_out15 <= XSIG591;
						i <= i + 1;
					WHEN 37 =>
						shift_out0 <= XSIG592;
						shift_out1 <= XSIG593;
						shift_out2 <= XSIG594;
						shift_out3 <= XSIG595;
						shift_out4 <= XSIG596;
						shift_out5 <= XSIG597;
						shift_out6 <= XSIG598;
						shift_out7 <= XSIG599;
						shift_out8 <= XSIG600;
						shift_out9 <= XSIG601;
						shift_out10 <= XSIG602;
						shift_out11 <= XSIG603;
						shift_out12 <= XSIG604;
						shift_out13 <= XSIG605;
						shift_out14 <= XSIG606;
						shift_out15 <= XSIG607;
						i <= i + 1;
					WHEN 38 =>
						shift_out0 <= XSIG608;
						shift_out1 <= XSIG609;
						shift_out2 <= XSIG610;
						shift_out3 <= XSIG611;
						shift_out4 <= XSIG612;
						shift_out5 <= XSIG613;
						shift_out6 <= XSIG614;
						shift_out7 <= XSIG615;
						shift_out8 <= XSIG616;
						shift_out9 <= XSIG617;
						shift_out10 <= XSIG618;
						shift_out11 <= XSIG619;
						shift_out12 <= XSIG620;
						shift_out13 <= XSIG621;
						shift_out14 <= XSIG622;
						shift_out15 <= XSIG623;
						i <= i + 1;
					WHEN 39 =>
						shift_out0 <= XSIG624;
						shift_out1 <= XSIG625;
						shift_out2 <= XSIG626;
						shift_out3 <= XSIG627;
						shift_out4 <= XSIG628;
						shift_out5 <= XSIG629;
						shift_out6 <= XSIG630;
						shift_out7 <= XSIG631;
						shift_out8 <= XSIG632;
						shift_out9 <= XSIG633;
						shift_out10 <= XSIG634;
						shift_out11 <= XSIG635;
						shift_out12 <= XSIG636;
						shift_out13 <= XSIG637;
						shift_out14 <= XSIG638;
						shift_out15 <= XSIG639;
						i <= i + 1;
					WHEN 40 =>
						shift_out0 <= XSIG640;
						shift_out1 <= XSIG641;
						shift_out2 <= XSIG642;
						shift_out3 <= XSIG643;
						shift_out4 <= XSIG644;
						shift_out5 <= XSIG645;
						shift_out6 <= XSIG646;
						shift_out7 <= XSIG647;
						shift_out8 <= XSIG648;
						shift_out9 <= XSIG649;
						shift_out10 <= XSIG650;
						shift_out11 <= XSIG651;
						shift_out12 <= XSIG652;
						shift_out13 <= XSIG653;
						shift_out14 <= XSIG654;
						shift_out15 <= XSIG655;
						i <= i + 1;
					WHEN 41 =>
						shift_out0 <= XSIG656;
						shift_out1 <= XSIG657;
						shift_out2 <= XSIG658;
						shift_out3 <= XSIG659;
						shift_out4 <= XSIG660;
						shift_out5 <= XSIG661;
						shift_out6 <= XSIG662;
						shift_out7 <= XSIG663;
						shift_out8 <= XSIG664;
						shift_out9 <= XSIG665;
						shift_out10 <= XSIG666;
						shift_out11 <= XSIG667;
						shift_out12 <= XSIG668;
						shift_out13 <= XSIG669;
						shift_out14 <= XSIG670;
						shift_out15 <= XSIG671;
						i <= i + 1;
					WHEN 42 =>
						shift_out0 <= XSIG672;
						shift_out1 <= XSIG673;
						shift_out2 <= XSIG674;
						shift_out3 <= XSIG675;
						shift_out4 <= XSIG676;
						shift_out5 <= XSIG677;
						shift_out6 <= XSIG678;
						shift_out7 <= XSIG679;
						shift_out8 <= XSIG680;
						shift_out9 <= XSIG681;
						shift_out10 <= XSIG682;
						shift_out11 <= XSIG683;
						shift_out12 <= XSIG684;
						shift_out13 <= XSIG685;
						shift_out14 <= XSIG686;
						shift_out15 <= XSIG687;
						i <= i + 1;
					WHEN 43 =>
						shift_out0 <= XSIG688;
						shift_out1 <= XSIG689;
						shift_out2 <= XSIG690;
						shift_out3 <= XSIG691;
						shift_out4 <= XSIG692;
						shift_out5 <= XSIG693;
						shift_out6 <= XSIG694;
						shift_out7 <= XSIG695;
						shift_out8 <= XSIG696;
						shift_out9 <= XSIG697;
						shift_out10 <= XSIG698;
						shift_out11 <= XSIG699;
						shift_out12 <= XSIG700;
						shift_out13 <= XSIG701;
						shift_out14 <= XSIG702;
						shift_out15 <= XSIG703;
						i <= i + 1;
					WHEN 44 =>
						shift_out0 <= XSIG704;
						shift_out1 <= XSIG705;
						shift_out2 <= XSIG706;
						shift_out3 <= XSIG707;
						shift_out4 <= XSIG708;
						shift_out5 <= XSIG709;
						shift_out6 <= XSIG710;
						shift_out7 <= XSIG711;
						shift_out8 <= XSIG712;
						shift_out9 <= XSIG713;
						shift_out10 <= XSIG714;
						shift_out11 <= XSIG715;
						shift_out12 <= XSIG716;
						shift_out13 <= XSIG717;
						shift_out14 <= XSIG718;
						shift_out15 <= XSIG719;
						i <= i + 1;
					WHEN 45 =>
						shift_out0 <= XSIG720;
						shift_out1 <= XSIG721;
						shift_out2 <= XSIG722;
						shift_out3 <= XSIG723;
						shift_out4 <= XSIG724;
						shift_out5 <= XSIG725;
						shift_out6 <= XSIG726;
						shift_out7 <= XSIG727;
						shift_out8 <= XSIG728;
						shift_out9 <= XSIG729;
						shift_out10 <= XSIG730;
						shift_out11 <= XSIG731;
						shift_out12 <= XSIG732;
						shift_out13 <= XSIG733;
						shift_out14 <= XSIG734;
						shift_out15 <= XSIG735;
						i <= i + 1;
					WHEN 46 =>
						shift_out0 <= XSIG736;
						shift_out1 <= XSIG737;
						shift_out2 <= XSIG738;
						shift_out3 <= XSIG739;
						shift_out4 <= XSIG740;
						shift_out5 <= XSIG741;
						shift_out6 <= XSIG742;
						shift_out7 <= XSIG743;
						shift_out8 <= XSIG744;
						shift_out9 <= XSIG745;
						shift_out10 <= XSIG746;
						shift_out11 <= XSIG747;
						shift_out12 <= XSIG748;
						shift_out13 <= XSIG749;
						shift_out14 <= XSIG750;
						shift_out15 <= XSIG751;
						i <= i + 1;
					WHEN 47 =>
						shift_out0 <= XSIG752;
						shift_out1 <= XSIG753;
						shift_out2 <= XSIG754;
						shift_out3 <= XSIG755;
						shift_out4 <= XSIG756;
						shift_out5 <= XSIG757;
						shift_out6 <= XSIG758;
						shift_out7 <= XSIG759;
						shift_out8 <= XSIG760;
						shift_out9 <= XSIG761;
						shift_out10 <= XSIG762;
						shift_out11 <= XSIG763;
						shift_out12 <= XSIG764;
						shift_out13 <= XSIG765;
						shift_out14 <= XSIG766;
						shift_out15 <= XSIG767;
						i <= i + 1;
					WHEN 48 =>
						shift_out0 <= XSIG768;
						shift_out1 <= XSIG769;
						shift_out2 <= XSIG770;
						shift_out3 <= XSIG771;
						shift_out4 <= XSIG772;
						shift_out5 <= XSIG773;
						shift_out6 <= XSIG774;
						shift_out7 <= XSIG775;
						shift_out8 <= XSIG776;
						shift_out9 <= XSIG777;
						shift_out10 <= XSIG778;
						shift_out11 <= XSIG779;
						shift_out12 <= XSIG780;
						shift_out13 <= XSIG781;
						shift_out14 <= XSIG782;
						shift_out15 <= XSIG783;
						i <= i + 1;
					WHEN 49 =>
						shift_out0 <= XSIG784;
						shift_out1 <= XSIG785;
						shift_out2 <= XSIG786;
						shift_out3 <= XSIG787;
						shift_out4 <= XSIG788;
						shift_out5 <= XSIG789;
						shift_out6 <= XSIG790;
						shift_out7 <= XSIG791;
						shift_out8 <= XSIG792;
						shift_out9 <= XSIG793;
						shift_out10 <= XSIG794;
						shift_out11 <= XSIG795;
						shift_out12 <= XSIG796;
						shift_out13 <= XSIG797;
						shift_out14 <= XSIG798;
						shift_out15 <= XSIG799;
						i <= i + 1;
					WHEN 50 =>
						shift_out0 <= XSIG800;
						shift_out1 <= XSIG801;
						shift_out2 <= XSIG802;
						shift_out3 <= XSIG803;
						shift_out4 <= XSIG804;
						shift_out5 <= XSIG805;
						shift_out6 <= XSIG806;
						shift_out7 <= XSIG807;
						shift_out8 <= XSIG808;
						shift_out9 <= XSIG809;
						shift_out10 <= XSIG810;
						shift_out11 <= XSIG811;
						shift_out12 <= XSIG812;
						shift_out13 <= XSIG813;
						shift_out14 <= XSIG814;
						shift_out15 <= XSIG815;
						i <= i + 1;
					WHEN 51 =>
						shift_out0 <= XSIG816;
						shift_out1 <= XSIG817;
						shift_out2 <= XSIG818;
						shift_out3 <= XSIG819;
						shift_out4 <= XSIG820;
						shift_out5 <= XSIG821;
						shift_out6 <= XSIG822;
						shift_out7 <= XSIG823;
						shift_out8 <= XSIG824;
						shift_out9 <= XSIG825;
						shift_out10 <= XSIG826;
						shift_out11 <= XSIG827;
						shift_out12 <= XSIG828;
						shift_out13 <= XSIG829;
						shift_out14 <= XSIG830;
						shift_out15 <= XSIG831;
						i <= i + 1;
					WHEN 52 =>
						shift_out0 <= XSIG832;
						shift_out1 <= XSIG833;
						shift_out2 <= XSIG834;
						shift_out3 <= XSIG835;
						shift_out4 <= XSIG836;
						shift_out5 <= XSIG837;
						shift_out6 <= XSIG838;
						shift_out7 <= XSIG839;
						shift_out8 <= XSIG840;
						shift_out9 <= XSIG841;
						shift_out10 <= XSIG842;
						shift_out11 <= XSIG843;
						shift_out12 <= XSIG844;
						shift_out13 <= XSIG845;
						shift_out14 <= XSIG846;
						shift_out15 <= XSIG847;
						i <= i + 1;
					WHEN 53 =>
						shift_out0 <= XSIG848;
						shift_out1 <= XSIG849;
						shift_out2 <= XSIG850;
						shift_out3 <= XSIG851;
						shift_out4 <= XSIG852;
						shift_out5 <= XSIG853;
						shift_out6 <= XSIG854;
						shift_out7 <= XSIG855;
						shift_out8 <= XSIG856;
						shift_out9 <= XSIG857;
						shift_out10 <= XSIG858;
						shift_out11 <= XSIG859;
						shift_out12 <= XSIG860;
						shift_out13 <= XSIG861;
						shift_out14 <= XSIG862;
						shift_out15 <= XSIG863;
						i <= i + 1;
					WHEN 54 =>
						shift_out0 <= XSIG864;
						shift_out1 <= XSIG865;
						shift_out2 <= XSIG866;
						shift_out3 <= XSIG867;
						shift_out4 <= XSIG868;
						shift_out5 <= XSIG869;
						shift_out6 <= XSIG870;
						shift_out7 <= XSIG871;
						shift_out8 <= XSIG872;
						shift_out9 <= XSIG873;
						shift_out10 <= XSIG874;
						shift_out11 <= XSIG875;
						shift_out12 <= XSIG876;
						shift_out13 <= XSIG877;
						shift_out14 <= XSIG878;
						shift_out15 <= XSIG879;
						i <= i + 1;
					WHEN 55 =>
						shift_out0 <= XSIG880;
						shift_out1 <= XSIG881;
						shift_out2 <= XSIG882;
						shift_out3 <= XSIG883;
						shift_out4 <= XSIG884;
						shift_out5 <= XSIG885;
						shift_out6 <= XSIG886;
						shift_out7 <= XSIG887;
						shift_out8 <= XSIG888;
						shift_out9 <= XSIG889;
						shift_out10 <= XSIG890;
						shift_out11 <= XSIG891;
						shift_out12 <= XSIG892;
						shift_out13 <= XSIG893;
						shift_out14 <= XSIG894;
						shift_out15 <= XSIG895;
						i <= i + 1;
					WHEN 56 =>
						shift_out0 <= XSIG896;
						shift_out1 <= XSIG897;
						shift_out2 <= XSIG898;
						shift_out3 <= XSIG899;
						shift_out4 <= XSIG900;
						shift_out5 <= XSIG901;
						shift_out6 <= XSIG902;
						shift_out7 <= XSIG903;
						shift_out8 <= XSIG904;
						shift_out9 <= XSIG905;
						shift_out10 <= XSIG906;
						shift_out11 <= XSIG907;
						shift_out12 <= XSIG908;
						shift_out13 <= XSIG909;
						shift_out14 <= XSIG910;
						shift_out15 <= XSIG911;
						i <= i + 1;
					WHEN 57 =>
						shift_out0 <= XSIG912;
						shift_out1 <= XSIG913;
						shift_out2 <= XSIG914;
						shift_out3 <= XSIG915;
						shift_out4 <= XSIG916;
						shift_out5 <= XSIG917;
						shift_out6 <= XSIG918;
						shift_out7 <= XSIG919;
						shift_out8 <= XSIG920;
						shift_out9 <= XSIG921;
						shift_out10 <= XSIG922;
						shift_out11 <= XSIG923;
						shift_out12 <= XSIG924;
						shift_out13 <= XSIG925;
						shift_out14 <= XSIG926;
						shift_out15 <= XSIG927;
						i <= i + 1;
					WHEN 58 =>
						shift_out0 <= XSIG928;
						shift_out1 <= XSIG929;
						shift_out2 <= XSIG930;
						shift_out3 <= XSIG931;
						shift_out4 <= XSIG932;
						shift_out5 <= XSIG933;
						shift_out6 <= XSIG934;
						shift_out7 <= XSIG935;
						shift_out8 <= XSIG936;
						shift_out9 <= XSIG937;
						shift_out10 <= XSIG938;
						shift_out11 <= XSIG939;
						shift_out12 <= XSIG940;
						shift_out13 <= XSIG941;
						shift_out14 <= XSIG942;
						shift_out15 <= XSIG943;
						i <= i + 1;
					WHEN 59 =>
						shift_out0 <= XSIG944;
						shift_out1 <= XSIG945;
						shift_out2 <= XSIG946;
						shift_out3 <= XSIG947;
						shift_out4 <= XSIG948;
						shift_out5 <= XSIG949;
						shift_out6 <= XSIG950;
						shift_out7 <= XSIG951;
						shift_out8 <= XSIG952;
						shift_out9 <= XSIG953;
						shift_out10 <= XSIG954;
						shift_out11 <= XSIG955;
						shift_out12 <= XSIG956;
						shift_out13 <= XSIG957;
						shift_out14 <= XSIG958;
						shift_out15 <= XSIG959;
						i <= i + 1;
					WHEN 60 =>
						shift_out0 <= XSIG960;
						shift_out1 <= XSIG961;
						shift_out2 <= XSIG962;
						shift_out3 <= XSIG963;
						shift_out4 <= XSIG964;
						shift_out5 <= XSIG965;
						shift_out6 <= XSIG966;
						shift_out7 <= XSIG967;
						shift_out8 <= XSIG968;
						shift_out9 <= XSIG969;
						shift_out10 <= XSIG970;
						shift_out11 <= XSIG971;
						shift_out12 <= XSIG972;
						shift_out13 <= XSIG973;
						shift_out14 <= XSIG974;
						shift_out15 <= XSIG975;
						i <= i + 1;
					WHEN 61 =>
						shift_out0 <= XSIG976;
						shift_out1 <= XSIG977;
						shift_out2 <= XSIG978;
						shift_out3 <= XSIG979;
						shift_out4 <= XSIG980;
						shift_out5 <= XSIG981;
						shift_out6 <= XSIG982;
						shift_out7 <= XSIG983;
						shift_out8 <= XSIG984;
						shift_out9 <= XSIG985;
						shift_out10 <= XSIG986;
						shift_out11 <= XSIG987;
						shift_out12 <= XSIG988;
						shift_out13 <= XSIG989;
						shift_out14 <= XSIG990;
						shift_out15 <= XSIG991;
						i <= i + 1;
					WHEN 62 =>
						shift_out0 <= XSIG992;
						shift_out1 <= XSIG993;
						shift_out2 <= XSIG994;
						shift_out3 <= XSIG995;
						shift_out4 <= XSIG996;
						shift_out5 <= XSIG997;
						shift_out6 <= XSIG998;
						shift_out7 <= XSIG999;
						shift_out8 <= XSIG1000;
						shift_out9 <= XSIG1001;
						shift_out10 <= XSIG1002;
						shift_out11 <= XSIG1003;
						shift_out12 <= XSIG1004;
						shift_out13 <= XSIG1005;
						shift_out14 <= XSIG1006;
						shift_out15 <= XSIG1007;
						i <= i + 1;
					WHEN 63 =>
						shift_out0 <= XSIG1008;
						shift_out1 <= XSIG1009;
						shift_out2 <= XSIG1010;
						shift_out3 <= XSIG1011;
						shift_out4 <= XSIG1012;
						shift_out5 <= XSIG1013;
						shift_out6 <= XSIG1014;
						shift_out7 <= XSIG1015;
						shift_out8 <= XSIG1016;
						shift_out9 <= XSIG1017;
						shift_out10 <= XSIG1018;
						shift_out11 <= XSIG1019;
						shift_out12 <= XSIG1020;
						shift_out13 <= XSIG1021;
						shift_out14 <= XSIG1022;
						shift_out15 <= XSIG1023;
						i <= i + 1;
					WHEN 64 =>
						shift_out0 <= XSIG1024;
						shift_out1 <= XSIG1025;
						shift_out2 <= XSIG1026;
						shift_out3 <= XSIG1027;
						shift_out4 <= XSIG1028;
						shift_out5 <= XSIG1029;
						shift_out6 <= XSIG1030;
						shift_out7 <= XSIG1031;
						shift_out8 <= XSIG1032;
						shift_out9 <= XSIG1033;
						shift_out10 <= XSIG1034;
						shift_out11 <= XSIG1035;
						shift_out12 <= XSIG1036;
						shift_out13 <= XSIG1037;
						shift_out14 <= XSIG1038;
						shift_out15 <= XSIG1039;
						i <= i + 1;
					WHEN 65 =>
						shift_out0 <= XSIG1040;
						shift_out1 <= XSIG1041;
						shift_out2 <= XSIG1042;
						shift_out3 <= XSIG1043;
						shift_out4 <= XSIG1044;
						shift_out5 <= XSIG1045;
						shift_out6 <= XSIG1046;
						shift_out7 <= XSIG1047;
						shift_out8 <= XSIG1048;
						shift_out9 <= XSIG1049;
						shift_out10 <= XSIG1050;
						shift_out11 <= XSIG1051;
						shift_out12 <= XSIG1052;
						shift_out13 <= XSIG1053;
						shift_out14 <= XSIG1054;
						shift_out15 <= XSIG1055;
						i <= i + 1;
					WHEN 66 =>
						shift_out0 <= XSIG1056;
						shift_out1 <= XSIG1057;
						shift_out2 <= XSIG1058;
						shift_out3 <= XSIG1059;
						shift_out4 <= XSIG1060;
						shift_out5 <= XSIG1061;
						shift_out6 <= XSIG1062;
						shift_out7 <= XSIG1063;
						shift_out8 <= XSIG1064;
						shift_out9 <= XSIG1065;
						shift_out10 <= XSIG1066;
						shift_out11 <= XSIG1067;
						shift_out12 <= XSIG1068;
						shift_out13 <= XSIG1069;
						shift_out14 <= XSIG1070;
						shift_out15 <= XSIG1071;
						i <= i + 1;
					WHEN 67 =>
						shift_out0 <= XSIG1072;
						shift_out1 <= XSIG1073;
						shift_out2 <= XSIG1074;
						shift_out3 <= XSIG1075;
						shift_out4 <= XSIG1076;
						shift_out5 <= XSIG1077;
						shift_out6 <= XSIG1078;
						shift_out7 <= XSIG1079;
						shift_out8 <= XSIG1080;
						shift_out9 <= XSIG1081;
						shift_out10 <= XSIG1082;
						shift_out11 <= XSIG1083;
						shift_out12 <= XSIG1084;
						shift_out13 <= XSIG1085;
						shift_out14 <= XSIG1086;
						shift_out15 <= XSIG1087;
						i <= i + 1;
					WHEN 68 =>
						shift_out0 <= XSIG1088;
						shift_out1 <= XSIG1089;
						shift_out2 <= XSIG1090;
						shift_out3 <= XSIG1091;
						shift_out4 <= XSIG1092;
						shift_out5 <= XSIG1093;
						shift_out6 <= XSIG1094;
						shift_out7 <= XSIG1095;
						shift_out8 <= XSIG1096;
						shift_out9 <= XSIG1097;
						shift_out10 <= XSIG1098;
						shift_out11 <= XSIG1099;
						shift_out12 <= XSIG1100;
						shift_out13 <= XSIG1101;
						shift_out14 <= XSIG1102;
						shift_out15 <= XSIG1103;
						i <= i + 1;
					WHEN 69 =>
						shift_out0 <= XSIG1104;
						shift_out1 <= XSIG1105;
						shift_out2 <= XSIG1106;
						shift_out3 <= XSIG1107;
						shift_out4 <= XSIG1108;
						shift_out5 <= XSIG1109;
						shift_out6 <= XSIG1110;
						shift_out7 <= XSIG1111;
						shift_out8 <= XSIG1112;
						shift_out9 <= XSIG1113;
						shift_out10 <= XSIG1114;
						shift_out11 <= XSIG1115;
						shift_out12 <= XSIG1116;
						shift_out13 <= XSIG1117;
						shift_out14 <= XSIG1118;
						shift_out15 <= XSIG1119;
						i <= i + 1;
					WHEN 70 =>
						shift_out0 <= XSIG1120;
						shift_out1 <= XSIG1121;
						shift_out2 <= XSIG1122;
						shift_out3 <= XSIG1123;
						shift_out4 <= XSIG1124;
						shift_out5 <= XSIG1125;
						shift_out6 <= XSIG1126;
						shift_out7 <= XSIG1127;
						shift_out8 <= XSIG1128;
						shift_out9 <= XSIG1129;
						shift_out10 <= XSIG1130;
						shift_out11 <= XSIG1131;
						shift_out12 <= XSIG1132;
						shift_out13 <= XSIG1133;
						shift_out14 <= XSIG1134;
						shift_out15 <= XSIG1135;
						i <= i + 1;
					WHEN 71 =>
						shift_out0 <= XSIG1136;
						shift_out1 <= XSIG1137;
						shift_out2 <= XSIG1138;
						shift_out3 <= XSIG1139;
						shift_out4 <= XSIG1140;
						shift_out5 <= XSIG1141;
						shift_out6 <= XSIG1142;
						shift_out7 <= XSIG1143;
						shift_out8 <= XSIG1144;
						shift_out9 <= XSIG1145;
						shift_out10 <= XSIG1146;
						shift_out11 <= XSIG1147;
						shift_out12 <= XSIG1148;
						shift_out13 <= XSIG1149;
						shift_out14 <= XSIG1150;
						shift_out15 <= XSIG1151;
						i <= i + 1;
					WHEN 72 =>
						shift_out0 <= XSIG1152;
						shift_out1 <= XSIG1153;
						shift_out2 <= XSIG1154;
						shift_out3 <= XSIG1155;
						shift_out4 <= XSIG1156;
						shift_out5 <= XSIG1157;
						shift_out6 <= XSIG1158;
						shift_out7 <= XSIG1159;
						shift_out8 <= XSIG1160;
						shift_out9 <= XSIG1161;
						shift_out10 <= XSIG1162;
						shift_out11 <= XSIG1163;
						shift_out12 <= XSIG1164;
						shift_out13 <= XSIG1165;
						shift_out14 <= XSIG1166;
						shift_out15 <= XSIG1167;
						i <= i + 1;
					WHEN 73 =>
						shift_out0 <= XSIG1168;
						shift_out1 <= XSIG1169;
						shift_out2 <= XSIG1170;
						shift_out3 <= XSIG1171;
						shift_out4 <= XSIG1172;
						shift_out5 <= XSIG1173;
						shift_out6 <= XSIG1174;
						shift_out7 <= XSIG1175;
						shift_out8 <= XSIG1176;
						shift_out9 <= XSIG1177;
						shift_out10 <= XSIG1178;
						shift_out11 <= XSIG1179;
						shift_out12 <= XSIG1180;
						shift_out13 <= XSIG1181;
						shift_out14 <= XSIG1182;
						shift_out15 <= XSIG1183;
						i <= i + 1;
					WHEN 74 =>
						shift_out0 <= XSIG1184;
						shift_out1 <= XSIG1185;
						shift_out2 <= XSIG1186;
						shift_out3 <= XSIG1187;
						shift_out4 <= XSIG1188;
						shift_out5 <= XSIG1189;
						shift_out6 <= XSIG1190;
						shift_out7 <= XSIG1191;
						shift_out8 <= XSIG1192;
						shift_out9 <= XSIG1193;
						shift_out10 <= XSIG1194;
						shift_out11 <= XSIG1195;
						shift_out12 <= XSIG1196;
						shift_out13 <= XSIG1197;
						shift_out14 <= XSIG1198;
						shift_out15 <= XSIG1199;
						i <= i + 1;
					WHEN 75 =>
						shift_out0 <= XSIG1200;
						shift_out1 <= XSIG1201;
						shift_out2 <= XSIG1202;
						shift_out3 <= XSIG1203;
						shift_out4 <= XSIG1204;
						shift_out5 <= XSIG1205;
						shift_out6 <= XSIG1206;
						shift_out7 <= XSIG1207;
						shift_out8 <= XSIG1208;
						shift_out9 <= XSIG1209;
						shift_out10 <= XSIG1210;
						shift_out11 <= XSIG1211;
						shift_out12 <= XSIG1212;
						shift_out13 <= XSIG1213;
						shift_out14 <= XSIG1214;
						shift_out15 <= XSIG1215;
						i <= i + 1;
					WHEN 76 =>
						shift_out0 <= XSIG1216;
						shift_out1 <= XSIG1217;
						shift_out2 <= XSIG1218;
						shift_out3 <= XSIG1219;
						shift_out4 <= XSIG1220;
						shift_out5 <= XSIG1221;
						shift_out6 <= XSIG1222;
						shift_out7 <= XSIG1223;
						shift_out8 <= XSIG1224;
						shift_out9 <= XSIG1225;
						shift_out10 <= XSIG1226;
						shift_out11 <= XSIG1227;
						shift_out12 <= XSIG1228;
						shift_out13 <= XSIG1229;
						shift_out14 <= XSIG1230;
						shift_out15 <= XSIG1231;
						i <= i + 1;
					WHEN 77 =>
						shift_out0 <= XSIG1232;
						shift_out1 <= XSIG1233;
						shift_out2 <= XSIG1234;
						shift_out3 <= XSIG1235;
						shift_out4 <= XSIG1236;
						shift_out5 <= XSIG1237;
						shift_out6 <= XSIG1238;
						shift_out7 <= XSIG1239;
						shift_out8 <= XSIG1240;
						shift_out9 <= XSIG1241;
						shift_out10 <= XSIG1242;
						shift_out11 <= XSIG1243;
						shift_out12 <= XSIG1244;
						shift_out13 <= XSIG1245;
						shift_out14 <= XSIG1246;
						shift_out15 <= XSIG1247;
						i <= i + 1;
					WHEN 78 =>
						shift_out0 <= XSIG1248;
						shift_out1 <= XSIG1249;
						shift_out2 <= XSIG1250;
						shift_out3 <= XSIG1251;
						shift_out4 <= XSIG1252;
						shift_out5 <= XSIG1253;
						shift_out6 <= XSIG1254;
						shift_out7 <= XSIG1255;
						shift_out8 <= XSIG1256;
						shift_out9 <= XSIG1257;
						shift_out10 <= XSIG1258;
						shift_out11 <= XSIG1259;
						shift_out12 <= XSIG1260;
						shift_out13 <= XSIG1261;
						shift_out14 <= XSIG1262;
						shift_out15 <= XSIG1263;
						i <= i + 1;
					WHEN 79 =>
						shift_out0 <= XSIG1264;
						shift_out1 <= XSIG1265;
						shift_out2 <= XSIG1266;
						shift_out3 <= XSIG1267;
						shift_out4 <= XSIG1268;
						shift_out5 <= XSIG1269;
						shift_out6 <= XSIG1270;
						shift_out7 <= XSIG1271;
						shift_out8 <= XSIG1272;
						shift_out9 <= XSIG1273;
						shift_out10 <= XSIG1274;
						shift_out11 <= XSIG1275;
						shift_out12 <= XSIG1276;
						shift_out13 <= XSIG1277;
						shift_out14 <= XSIG1278;
						shift_out15 <= XSIG1279;
						i <= i + 1;
					WHEN 80 =>
						shift_out0 <= XSIG1280;
						shift_out1 <= XSIG1281;
						shift_out2 <= XSIG1282;
						shift_out3 <= XSIG1283;
						shift_out4 <= XSIG1284;
						shift_out5 <= XSIG1285;
						shift_out6 <= XSIG1286;
						shift_out7 <= XSIG1287;
						shift_out8 <= XSIG1288;
						shift_out9 <= XSIG1289;
						shift_out10 <= XSIG1290;
						shift_out11 <= XSIG1291;
						shift_out12 <= XSIG1292;
						shift_out13 <= XSIG1293;
						shift_out14 <= XSIG1294;
						shift_out15 <= XSIG1295;
						i <= i + 1;
					WHEN 81 =>
						shift_out0 <= XSIG1296;
						shift_out1 <= XSIG1297;
						shift_out2 <= XSIG1298;
						shift_out3 <= XSIG1299;
						shift_out4 <= XSIG1300;
						shift_out5 <= XSIG1301;
						shift_out6 <= XSIG1302;
						shift_out7 <= XSIG1303;
						shift_out8 <= XSIG1304;
						shift_out9 <= XSIG1305;
						shift_out10 <= XSIG1306;
						shift_out11 <= XSIG1307;
						shift_out12 <= XSIG1308;
						shift_out13 <= XSIG1309;
						shift_out14 <= XSIG1310;
						shift_out15 <= XSIG1311;
						i <= i + 1;
					WHEN 82 =>
						shift_out0 <= XSIG1312;
						shift_out1 <= XSIG1313;
						shift_out2 <= XSIG1314;
						shift_out3 <= XSIG1315;
						shift_out4 <= XSIG1316;
						shift_out5 <= XSIG1317;
						shift_out6 <= XSIG1318;
						shift_out7 <= XSIG1319;
						shift_out8 <= XSIG1320;
						shift_out9 <= XSIG1321;
						shift_out10 <= XSIG1322;
						shift_out11 <= XSIG1323;
						shift_out12 <= XSIG1324;
						shift_out13 <= XSIG1325;
						shift_out14 <= XSIG1326;
						shift_out15 <= XSIG1327;
						i <= i + 1;
					WHEN 83 =>
						shift_out0 <= XSIG1328;
						shift_out1 <= XSIG1329;
						shift_out2 <= XSIG1330;
						shift_out3 <= XSIG1331;
						shift_out4 <= XSIG1332;
						shift_out5 <= XSIG1333;
						shift_out6 <= XSIG1334;
						shift_out7 <= XSIG1335;
						shift_out8 <= XSIG1336;
						shift_out9 <= XSIG1337;
						shift_out10 <= XSIG1338;
						shift_out11 <= XSIG1339;
						shift_out12 <= XSIG1340;
						shift_out13 <= XSIG1341;
						shift_out14 <= XSIG1342;
						shift_out15 <= XSIG1343;
						i <= i + 1;
					WHEN 84 =>
						shift_out0 <= XSIG1344;
						shift_out1 <= XSIG1345;
						shift_out2 <= XSIG1346;
						shift_out3 <= XSIG1347;
						shift_out4 <= XSIG1348;
						shift_out5 <= XSIG1349;
						shift_out6 <= XSIG1350;
						shift_out7 <= XSIG1351;
						shift_out8 <= XSIG1352;
						shift_out9 <= XSIG1353;
						shift_out10 <= XSIG1354;
						shift_out11 <= XSIG1355;
						shift_out12 <= XSIG1356;
						shift_out13 <= XSIG1357;
						shift_out14 <= XSIG1358;
						shift_out15 <= XSIG1359;
						i <= i + 1;
					WHEN 85 =>
						shift_out0 <= XSIG1360;
						shift_out1 <= XSIG1361;
						shift_out2 <= XSIG1362;
						shift_out3 <= XSIG1363;
						shift_out4 <= XSIG1364;
						shift_out5 <= XSIG1365;
						shift_out6 <= XSIG1366;
						shift_out7 <= XSIG1367;
						shift_out8 <= XSIG1368;
						shift_out9 <= XSIG1369;
						shift_out10 <= XSIG1370;
						shift_out11 <= XSIG1371;
						shift_out12 <= XSIG1372;
						shift_out13 <= XSIG1373;
						shift_out14 <= XSIG1374;
						shift_out15 <= XSIG1375;
						i <= i + 1;
					WHEN 86 =>
						shift_out0 <= XSIG1376;
						shift_out1 <= XSIG1377;
						shift_out2 <= XSIG1378;
						shift_out3 <= XSIG1379;
						shift_out4 <= XSIG1380;
						shift_out5 <= XSIG1381;
						shift_out6 <= XSIG1382;
						shift_out7 <= XSIG1383;
						shift_out8 <= XSIG1384;
						shift_out9 <= XSIG1385;
						shift_out10 <= XSIG1386;
						shift_out11 <= XSIG1387;
						shift_out12 <= XSIG1388;
						shift_out13 <= XSIG1389;
						shift_out14 <= XSIG1390;
						shift_out15 <= XSIG1391;
						i <= i + 1;
					WHEN 87 =>
						shift_out0 <= XSIG1392;
						shift_out1 <= XSIG1393;
						shift_out2 <= XSIG1394;
						shift_out3 <= XSIG1395;
						shift_out4 <= XSIG1396;
						shift_out5 <= XSIG1397;
						shift_out6 <= XSIG1398;
						shift_out7 <= XSIG1399;
						shift_out8 <= XSIG1400;
						shift_out9 <= XSIG1401;
						shift_out10 <= XSIG1402;
						shift_out11 <= XSIG1403;
						shift_out12 <= XSIG1404;
						shift_out13 <= XSIG1405;
						shift_out14 <= XSIG1406;
						shift_out15 <= XSIG1407;
						i <= i + 1;
					WHEN 88 =>
						shift_out0 <= XSIG1408;
						shift_out1 <= XSIG1409;
						shift_out2 <= XSIG1410;
						shift_out3 <= XSIG1411;
						shift_out4 <= XSIG1412;
						shift_out5 <= XSIG1413;
						shift_out6 <= XSIG1414;
						shift_out7 <= XSIG1415;
						shift_out8 <= XSIG1416;
						shift_out9 <= XSIG1417;
						shift_out10 <= XSIG1418;
						shift_out11 <= XSIG1419;
						shift_out12 <= XSIG1420;
						shift_out13 <= XSIG1421;
						shift_out14 <= XSIG1422;
						shift_out15 <= XSIG1423;
						i <= i + 1;
					WHEN 89 =>
						shift_out0 <= XSIG1424;
						shift_out1 <= XSIG1425;
						shift_out2 <= XSIG1426;
						shift_out3 <= XSIG1427;
						shift_out4 <= XSIG1428;
						shift_out5 <= XSIG1429;
						shift_out6 <= XSIG1430;
						shift_out7 <= XSIG1431;
						shift_out8 <= XSIG1432;
						shift_out9 <= XSIG1433;
						shift_out10 <= XSIG1434;
						shift_out11 <= XSIG1435;
						shift_out12 <= XSIG1436;
						shift_out13 <= XSIG1437;
						shift_out14 <= XSIG1438;
						shift_out15 <= XSIG1439;
						i <= i + 1;
					WHEN 90 =>
						shift_out0 <= XSIG1440;
						shift_out1 <= XSIG1441;
						shift_out2 <= XSIG1442;
						shift_out3 <= XSIG1443;
						shift_out4 <= XSIG1444;
						shift_out5 <= XSIG1445;
						shift_out6 <= XSIG1446;
						shift_out7 <= XSIG1447;
						shift_out8 <= XSIG1448;
						shift_out9 <= XSIG1449;
						shift_out10 <= XSIG1450;
						shift_out11 <= XSIG1451;
						shift_out12 <= XSIG1452;
						shift_out13 <= XSIG1453;
						shift_out14 <= XSIG1454;
						shift_out15 <= XSIG1455;
						i <= i + 1;
					WHEN 91 =>
						shift_out0 <= XSIG1456;
						shift_out1 <= XSIG1457;
						shift_out2 <= XSIG1458;
						shift_out3 <= XSIG1459;
						shift_out4 <= XSIG1460;
						shift_out5 <= XSIG1461;
						shift_out6 <= XSIG1462;
						shift_out7 <= XSIG1463;
						shift_out8 <= XSIG1464;
						shift_out9 <= XSIG1465;
						shift_out10 <= XSIG1466;
						shift_out11 <= XSIG1467;
						shift_out12 <= XSIG1468;
						shift_out13 <= XSIG1469;
						shift_out14 <= XSIG1470;
						shift_out15 <= XSIG1471;
						i <= i + 1;
					WHEN 92 =>
						shift_out0 <= XSIG1472;
						shift_out1 <= XSIG1473;
						shift_out2 <= XSIG1474;
						shift_out3 <= XSIG1475;
						shift_out4 <= XSIG1476;
						shift_out5 <= XSIG1477;
						shift_out6 <= XSIG1478;
						shift_out7 <= XSIG1479;
						shift_out8 <= XSIG1480;
						shift_out9 <= XSIG1481;
						shift_out10 <= XSIG1482;
						shift_out11 <= XSIG1483;
						shift_out12 <= XSIG1484;
						shift_out13 <= XSIG1485;
						shift_out14 <= XSIG1486;
						shift_out15 <= XSIG1487;
						i <= i + 1;
					WHEN 93 =>
						shift_out0 <= XSIG1488;
						shift_out1 <= XSIG1489;
						shift_out2 <= XSIG1490;
						shift_out3 <= XSIG1491;
						shift_out4 <= XSIG1492;
						shift_out5 <= XSIG1493;
						shift_out6 <= XSIG1494;
						shift_out7 <= XSIG1495;
						shift_out8 <= XSIG1496;
						shift_out9 <= XSIG1497;
						shift_out10 <= XSIG1498;
						shift_out11 <= XSIG1499;
						shift_out12 <= XSIG1500;
						shift_out13 <= XSIG1501;
						shift_out14 <= XSIG1502;
						shift_out15 <= XSIG1503;
						i <= i + 1;
					WHEN 94 =>
						shift_out0 <= XSIG1504;
						shift_out1 <= XSIG1505;
						shift_out2 <= XSIG1506;
						shift_out3 <= XSIG1507;
						shift_out4 <= XSIG1508;
						shift_out5 <= XSIG1509;
						shift_out6 <= XSIG1510;
						shift_out7 <= XSIG1511;
						shift_out8 <= XSIG1512;
						shift_out9 <= XSIG1513;
						shift_out10 <= XSIG1514;
						shift_out11 <= XSIG1515;
						shift_out12 <= XSIG1516;
						shift_out13 <= XSIG1517;
						shift_out14 <= XSIG1518;
						shift_out15 <= XSIG1519;
						i <= i + 1;
					WHEN 95 =>
						shift_out0 <= XSIG1520;
						shift_out1 <= XSIG1521;
						shift_out2 <= XSIG1522;
						shift_out3 <= XSIG1523;
						shift_out4 <= XSIG1524;
						shift_out5 <= XSIG1525;
						shift_out6 <= XSIG1526;
						shift_out7 <= XSIG1527;
						shift_out8 <= XSIG1528;
						shift_out9 <= XSIG1529;
						shift_out10 <= XSIG1530;
						shift_out11 <= XSIG1531;
						shift_out12 <= XSIG1532;
						shift_out13 <= XSIG1533;
						shift_out14 <= XSIG1534;
						shift_out15 <= XSIG1535;
						i <= i + 1;
					WHEN 96 =>
						shift_out0 <= XSIG1536;
						shift_out1 <= XSIG1537;
						shift_out2 <= XSIG1538;
						shift_out3 <= XSIG1539;
						shift_out4 <= XSIG1540;
						shift_out5 <= XSIG1541;
						shift_out6 <= XSIG1542;
						shift_out7 <= XSIG1543;
						shift_out8 <= XSIG1544;
						shift_out9 <= XSIG1545;
						shift_out10 <= XSIG1546;
						shift_out11 <= XSIG1547;
						shift_out12 <= XSIG1548;
						shift_out13 <= XSIG1549;
						shift_out14 <= XSIG1550;
						shift_out15 <= XSIG1551;
						i <= i + 1;
					WHEN 97 =>
						shift_out0 <= XSIG1552;
						shift_out1 <= XSIG1553;
						shift_out2 <= XSIG1554;
						shift_out3 <= XSIG1555;
						shift_out4 <= XSIG1556;
						shift_out5 <= XSIG1557;
						shift_out6 <= XSIG1558;
						shift_out7 <= XSIG1559;
						shift_out8 <= XSIG1560;
						shift_out9 <= XSIG1561;
						shift_out10 <= XSIG1562;
						shift_out11 <= XSIG1563;
						shift_out12 <= XSIG1564;
						shift_out13 <= XSIG1565;
						shift_out14 <= XSIG1566;
						shift_out15 <= XSIG1567;
						i <= i + 1;
					WHEN 98 =>
						shift_out0 <= XSIG1568;
						shift_out1 <= XSIG1569;
						shift_out2 <= XSIG1570;
						shift_out3 <= XSIG1571;
						shift_out4 <= XSIG1572;
						shift_out5 <= XSIG1573;
						shift_out6 <= XSIG1574;
						shift_out7 <= XSIG1575;
						shift_out8 <= XSIG1576;
						shift_out9 <= XSIG1577;
						shift_out10 <= XSIG1578;
						shift_out11 <= XSIG1579;
						shift_out12 <= XSIG1580;
						shift_out13 <= XSIG1581;
						shift_out14 <= XSIG1582;
						shift_out15 <= XSIG1583;
						i <= i + 1;
					WHEN 99 =>
						shift_out0 <= XSIG1584;
						shift_out1 <= XSIG1585;
						shift_out2 <= XSIG1586;
						shift_out3 <= XSIG1587;
						shift_out4 <= XSIG1588;
						shift_out5 <= XSIG1589;
						shift_out6 <= XSIG1590;
						shift_out7 <= XSIG1591;
						shift_out8 <= XSIG1592;
						shift_out9 <= XSIG1593;
						shift_out10 <= XSIG1594;
						shift_out11 <= XSIG1595;
						shift_out12 <= XSIG1596;
						shift_out13 <= XSIG1597;
						shift_out14 <= XSIG1598;
						shift_out15 <= XSIG1599;
						i <= i + 1;
					WHEN 100 =>
						shift_out0 <= XSIG1600;
						shift_out1 <= XSIG1601;
						shift_out2 <= XSIG1602;
						shift_out3 <= XSIG1603;
						shift_out4 <= XSIG1604;
						shift_out5 <= XSIG1605;
						shift_out6 <= XSIG1606;
						shift_out7 <= XSIG1607;
						shift_out8 <= XSIG1608;
						shift_out9 <= XSIG1609;
						shift_out10 <= XSIG1610;
						shift_out11 <= XSIG1611;
						shift_out12 <= XSIG1612;
						shift_out13 <= XSIG1613;
						shift_out14 <= XSIG1614;
						shift_out15 <= XSIG1615;
						i <= i + 1;
					WHEN 101 =>
						shift_out0 <= XSIG1616;
						shift_out1 <= XSIG1617;
						shift_out2 <= XSIG1618;
						shift_out3 <= XSIG1619;
						shift_out4 <= XSIG1620;
						shift_out5 <= XSIG1621;
						shift_out6 <= XSIG1622;
						shift_out7 <= XSIG1623;
						shift_out8 <= XSIG1624;
						shift_out9 <= XSIG1625;
						shift_out10 <= XSIG1626;
						shift_out11 <= XSIG1627;
						shift_out12 <= XSIG1628;
						shift_out13 <= XSIG1629;
						shift_out14 <= XSIG1630;
						shift_out15 <= XSIG1631;
						i <= i + 1;
					WHEN 102 =>
						shift_out0 <= XSIG1632;
						shift_out1 <= XSIG1633;
						shift_out2 <= XSIG1634;
						shift_out3 <= XSIG1635;
						shift_out4 <= XSIG1636;
						shift_out5 <= XSIG1637;
						shift_out6 <= XSIG1638;
						shift_out7 <= XSIG1639;
						shift_out8 <= XSIG1640;
						shift_out9 <= XSIG1641;
						shift_out10 <= XSIG1642;
						shift_out11 <= XSIG1643;
						shift_out12 <= XSIG1644;
						shift_out13 <= XSIG1645;
						shift_out14 <= XSIG1646;
						shift_out15 <= XSIG1647;
						i <= i + 1;
					WHEN 103 =>
						shift_out0 <= XSIG1648;
						shift_out1 <= XSIG1649;
						shift_out2 <= XSIG1650;
						shift_out3 <= XSIG1651;
						shift_out4 <= XSIG1652;
						shift_out5 <= XSIG1653;
						shift_out6 <= XSIG1654;
						shift_out7 <= XSIG1655;
						shift_out8 <= XSIG1656;
						shift_out9 <= XSIG1657;
						shift_out10 <= XSIG1658;
						shift_out11 <= XSIG1659;
						shift_out12 <= XSIG1660;
						shift_out13 <= XSIG1661;
						shift_out14 <= XSIG1662;
						shift_out15 <= XSIG1663;
						i <= i + 1;
					WHEN 104 =>
						shift_out0 <= XSIG1664;
						shift_out1 <= XSIG1665;
						shift_out2 <= XSIG1666;
						shift_out3 <= XSIG1667;
						shift_out4 <= XSIG1668;
						shift_out5 <= XSIG1669;
						shift_out6 <= XSIG1670;
						shift_out7 <= XSIG1671;
						shift_out8 <= XSIG1672;
						shift_out9 <= XSIG1673;
						shift_out10 <= XSIG1674;
						shift_out11 <= XSIG1675;
						shift_out12 <= XSIG1676;
						shift_out13 <= XSIG1677;
						shift_out14 <= XSIG1678;
						shift_out15 <= XSIG1679;
						i <= i + 1;
					WHEN 105 =>
						shift_out0 <= XSIG1680;
						shift_out1 <= XSIG1681;
						shift_out2 <= XSIG1682;
						shift_out3 <= XSIG1683;
						shift_out4 <= XSIG1684;
						shift_out5 <= XSIG1685;
						shift_out6 <= XSIG1686;
						shift_out7 <= XSIG1687;
						shift_out8 <= XSIG1688;
						shift_out9 <= XSIG1689;
						shift_out10 <= XSIG1690;
						shift_out11 <= XSIG1691;
						shift_out12 <= XSIG1692;
						shift_out13 <= XSIG1693;
						shift_out14 <= XSIG1694;
						shift_out15 <= XSIG1695;
						i <= i + 1;
					WHEN 106 =>
						shift_out0 <= XSIG1696;
						shift_out1 <= XSIG1697;
						shift_out2 <= XSIG1698;
						shift_out3 <= XSIG1699;
						shift_out4 <= XSIG1700;
						shift_out5 <= XSIG1701;
						shift_out6 <= XSIG1702;
						shift_out7 <= XSIG1703;
						shift_out8 <= XSIG1704;
						shift_out9 <= XSIG1705;
						shift_out10 <= XSIG1706;
						shift_out11 <= XSIG1707;
						shift_out12 <= XSIG1708;
						shift_out13 <= XSIG1709;
						shift_out14 <= XSIG1710;
						shift_out15 <= XSIG1711;
						i <= i + 1;
					WHEN 107 =>
						shift_out0 <= XSIG1712;
						shift_out1 <= XSIG1713;
						shift_out2 <= XSIG1714;
						shift_out3 <= XSIG1715;
						shift_out4 <= XSIG1716;
						shift_out5 <= XSIG1717;
						shift_out6 <= XSIG1718;
						shift_out7 <= XSIG1719;
						shift_out8 <= XSIG1720;
						shift_out9 <= XSIG1721;
						shift_out10 <= XSIG1722;
						shift_out11 <= XSIG1723;
						shift_out12 <= XSIG1724;
						shift_out13 <= XSIG1725;
						shift_out14 <= XSIG1726;
						shift_out15 <= XSIG1727;
						i <= i + 1;
					WHEN 108 =>
						shift_out0 <= XSIG1728;
						shift_out1 <= XSIG1729;
						shift_out2 <= XSIG1730;
						shift_out3 <= XSIG1731;
						shift_out4 <= XSIG1732;
						shift_out5 <= XSIG1733;
						shift_out6 <= XSIG1734;
						shift_out7 <= XSIG1735;
						shift_out8 <= XSIG1736;
						shift_out9 <= XSIG1737;
						shift_out10 <= XSIG1738;
						shift_out11 <= XSIG1739;
						shift_out12 <= XSIG1740;
						shift_out13 <= XSIG1741;
						shift_out14 <= XSIG1742;
						shift_out15 <= XSIG1743;
						i <= i + 1;
					WHEN 109 =>
						shift_out0 <= XSIG1744;
						shift_out1 <= XSIG1745;
						shift_out2 <= XSIG1746;
						shift_out3 <= XSIG1747;
						shift_out4 <= XSIG1748;
						shift_out5 <= XSIG1749;
						shift_out6 <= XSIG1750;
						shift_out7 <= XSIG1751;
						shift_out8 <= XSIG1752;
						shift_out9 <= XSIG1753;
						shift_out10 <= XSIG1754;
						shift_out11 <= XSIG1755;
						shift_out12 <= XSIG1756;
						shift_out13 <= XSIG1757;
						shift_out14 <= XSIG1758;
						shift_out15 <= XSIG1759;
						i <= i + 1;
					WHEN 110 =>
						shift_out0 <= XSIG1760;
						shift_out1 <= XSIG1761;
						shift_out2 <= XSIG1762;
						shift_out3 <= XSIG1763;
						shift_out4 <= XSIG1764;
						shift_out5 <= XSIG1765;
						shift_out6 <= XSIG1766;
						shift_out7 <= XSIG1767;
						shift_out8 <= XSIG1768;
						shift_out9 <= XSIG1769;
						shift_out10 <= XSIG1770;
						shift_out11 <= XSIG1771;
						shift_out12 <= XSIG1772;
						shift_out13 <= XSIG1773;
						shift_out14 <= XSIG1774;
						shift_out15 <= XSIG1775;
						i <= i + 1;
					WHEN 111 =>
						shift_out0 <= XSIG1776;
						shift_out1 <= XSIG1777;
						shift_out2 <= XSIG1778;
						shift_out3 <= XSIG1779;
						shift_out4 <= XSIG1780;
						shift_out5 <= XSIG1781;
						shift_out6 <= XSIG1782;
						shift_out7 <= XSIG1783;
						shift_out8 <= XSIG1784;
						shift_out9 <= XSIG1785;
						shift_out10 <= XSIG1786;
						shift_out11 <= XSIG1787;
						shift_out12 <= XSIG1788;
						shift_out13 <= XSIG1789;
						shift_out14 <= XSIG1790;
						shift_out15 <= XSIG1791;
						i <= i + 1;
					WHEN 112 =>
						shift_out0 <= XSIG1792;
						shift_out1 <= XSIG1793;
						shift_out2 <= XSIG1794;
						shift_out3 <= XSIG1795;
						shift_out4 <= XSIG1796;
						shift_out5 <= XSIG1797;
						shift_out6 <= XSIG1798;
						shift_out7 <= XSIG1799;
						shift_out8 <= XSIG1800;
						shift_out9 <= XSIG1801;
						shift_out10 <= XSIG1802;
						shift_out11 <= XSIG1803;
						shift_out12 <= XSIG1804;
						shift_out13 <= XSIG1805;
						shift_out14 <= XSIG1806;
						shift_out15 <= XSIG1807;
						i <= i + 1;
					WHEN 113 =>
						shift_out0 <= XSIG1808;
						shift_out1 <= XSIG1809;
						shift_out2 <= XSIG1810;
						shift_out3 <= XSIG1811;
						shift_out4 <= XSIG1812;
						shift_out5 <= XSIG1813;
						shift_out6 <= XSIG1814;
						shift_out7 <= XSIG1815;
						shift_out8 <= XSIG1816;
						shift_out9 <= XSIG1817;
						shift_out10 <= XSIG1818;
						shift_out11 <= XSIG1819;
						shift_out12 <= XSIG1820;
						shift_out13 <= XSIG1821;
						shift_out14 <= XSIG1822;
						shift_out15 <= XSIG1823;
						i <= i + 1;
					WHEN 114 =>
						shift_out0 <= XSIG1824;
						shift_out1 <= XSIG1825;
						shift_out2 <= XSIG1826;
						shift_out3 <= XSIG1827;
						shift_out4 <= XSIG1828;
						shift_out5 <= XSIG1829;
						shift_out6 <= XSIG1830;
						shift_out7 <= XSIG1831;
						shift_out8 <= XSIG1832;
						shift_out9 <= XSIG1833;
						shift_out10 <= XSIG1834;
						shift_out11 <= XSIG1835;
						shift_out12 <= XSIG1836;
						shift_out13 <= XSIG1837;
						shift_out14 <= XSIG1838;
						shift_out15 <= XSIG1839;
						i <= i + 1;
					WHEN 115 =>
						shift_out0 <= XSIG1840;
						shift_out1 <= XSIG1841;
						shift_out2 <= XSIG1842;
						shift_out3 <= XSIG1843;
						shift_out4 <= XSIG1844;
						shift_out5 <= XSIG1845;
						shift_out6 <= XSIG1846;
						shift_out7 <= XSIG1847;
						shift_out8 <= XSIG1848;
						shift_out9 <= XSIG1849;
						shift_out10 <= XSIG1850;
						shift_out11 <= XSIG1851;
						shift_out12 <= XSIG1852;
						shift_out13 <= XSIG1853;
						shift_out14 <= XSIG1854;
						shift_out15 <= XSIG1855;
						i <= i + 1;
					WHEN 116 =>
						shift_out0 <= XSIG1856;
						shift_out1 <= XSIG1857;
						shift_out2 <= XSIG1858;
						shift_out3 <= XSIG1859;
						shift_out4 <= XSIG1860;
						shift_out5 <= XSIG1861;
						shift_out6 <= XSIG1862;
						shift_out7 <= XSIG1863;
						shift_out8 <= XSIG1864;
						shift_out9 <= XSIG1865;
						shift_out10 <= XSIG1866;
						shift_out11 <= XSIG1867;
						shift_out12 <= XSIG1868;
						shift_out13 <= XSIG1869;
						shift_out14 <= XSIG1870;
						shift_out15 <= XSIG1871;
						i <= i + 1;
					WHEN 117 =>
						shift_out0 <= XSIG1872;
						shift_out1 <= XSIG1873;
						shift_out2 <= XSIG1874;
						shift_out3 <= XSIG1875;
						shift_out4 <= XSIG1876;
						shift_out5 <= XSIG1877;
						shift_out6 <= XSIG1878;
						shift_out7 <= XSIG1879;
						shift_out8 <= XSIG1880;
						shift_out9 <= XSIG1881;
						shift_out10 <= XSIG1882;
						shift_out11 <= XSIG1883;
						shift_out12 <= XSIG1884;
						shift_out13 <= XSIG1885;
						shift_out14 <= XSIG1886;
						shift_out15 <= XSIG1887;
						i <= i + 1;
					WHEN 118 =>
						shift_out0 <= XSIG1888;
						shift_out1 <= XSIG1889;
						shift_out2 <= XSIG1890;
						shift_out3 <= XSIG1891;
						shift_out4 <= XSIG1892;
						shift_out5 <= XSIG1893;
						shift_out6 <= XSIG1894;
						shift_out7 <= XSIG1895;
						shift_out8 <= XSIG1896;
						shift_out9 <= XSIG1897;
						shift_out10 <= XSIG1898;
						shift_out11 <= XSIG1899;
						shift_out12 <= XSIG1900;
						shift_out13 <= XSIG1901;
						shift_out14 <= XSIG1902;
						shift_out15 <= XSIG1903;
						i <= i + 1;
					WHEN 119 =>
						shift_out0 <= XSIG1904;
						shift_out1 <= XSIG1905;
						shift_out2 <= XSIG1906;
						shift_out3 <= XSIG1907;
						shift_out4 <= XSIG1908;
						shift_out5 <= XSIG1909;
						shift_out6 <= XSIG1910;
						shift_out7 <= XSIG1911;
						shift_out8 <= XSIG1912;
						shift_out9 <= XSIG1913;
						shift_out10 <= XSIG1914;
						shift_out11 <= XSIG1915;
						shift_out12 <= XSIG1916;
						shift_out13 <= XSIG1917;
						shift_out14 <= XSIG1918;
						shift_out15 <= XSIG1919;
						i <= i + 1;
					WHEN 120 =>
						shift_out0 <= XSIG1920;
						shift_out1 <= XSIG1921;
						shift_out2 <= XSIG1922;
						shift_out3 <= XSIG1923;
						shift_out4 <= XSIG1924;
						shift_out5 <= XSIG1925;
						shift_out6 <= XSIG1926;
						shift_out7 <= XSIG1927;
						shift_out8 <= XSIG1928;
						shift_out9 <= XSIG1929;
						shift_out10 <= XSIG1930;
						shift_out11 <= XSIG1931;
						shift_out12 <= XSIG1932;
						shift_out13 <= XSIG1933;
						shift_out14 <= XSIG1934;
						shift_out15 <= XSIG1935;
						i <= i + 1;
					WHEN 121 =>
						shift_out0 <= XSIG1936;
						shift_out1 <= XSIG1937;
						shift_out2 <= XSIG1938;
						shift_out3 <= XSIG1939;
						shift_out4 <= XSIG1940;
						shift_out5 <= XSIG1941;
						shift_out6 <= XSIG1942;
						shift_out7 <= XSIG1943;
						shift_out8 <= XSIG1944;
						shift_out9 <= XSIG1945;
						shift_out10 <= XSIG1946;
						shift_out11 <= XSIG1947;
						shift_out12 <= XSIG1948;
						shift_out13 <= XSIG1949;
						shift_out14 <= XSIG1950;
						shift_out15 <= XSIG1951;
						i <= i + 1;
					WHEN 122 =>
						shift_out0 <= XSIG1952;
						shift_out1 <= XSIG1953;
						shift_out2 <= XSIG1954;
						shift_out3 <= XSIG1955;
						shift_out4 <= XSIG1956;
						shift_out5 <= XSIG1957;
						shift_out6 <= XSIG1958;
						shift_out7 <= XSIG1959;
						shift_out8 <= XSIG1960;
						shift_out9 <= XSIG1961;
						shift_out10 <= XSIG1962;
						shift_out11 <= XSIG1963;
						shift_out12 <= XSIG1964;
						shift_out13 <= XSIG1965;
						shift_out14 <= XSIG1966;
						shift_out15 <= XSIG1967;
						i <= i + 1;
					WHEN 123 =>
						shift_out0 <= XSIG1968;
						shift_out1 <= XSIG1969;
						shift_out2 <= XSIG1970;
						shift_out3 <= XSIG1971;
						shift_out4 <= XSIG1972;
						shift_out5 <= XSIG1973;
						shift_out6 <= XSIG1974;
						shift_out7 <= XSIG1975;
						shift_out8 <= XSIG1976;
						shift_out9 <= XSIG1977;
						shift_out10 <= XSIG1978;
						shift_out11 <= XSIG1979;
						shift_out12 <= XSIG1980;
						shift_out13 <= XSIG1981;
						shift_out14 <= XSIG1982;
						shift_out15 <= XSIG1983;
						i <= i + 1;
					WHEN 124 =>
						shift_out0 <= XSIG1984;
						shift_out1 <= XSIG1985;
						shift_out2 <= XSIG1986;
						shift_out3 <= XSIG1987;
						shift_out4 <= XSIG1988;
						shift_out5 <= XSIG1989;
						shift_out6 <= XSIG1990;
						shift_out7 <= XSIG1991;
						shift_out8 <= XSIG1992;
						shift_out9 <= XSIG1993;
						shift_out10 <= XSIG1994;
						shift_out11 <= XSIG1995;
						shift_out12 <= XSIG1996;
						shift_out13 <= XSIG1997;
						shift_out14 <= XSIG1998;
						shift_out15 <= XSIG1999;
						i <= i + 1;
					WHEN 125 =>
						shift_out0 <= XSIG2000;
						shift_out1 <= XSIG2001;
						shift_out2 <= XSIG2002;
						shift_out3 <= XSIG2003;
						shift_out4 <= XSIG2004;
						shift_out5 <= XSIG2005;
						shift_out6 <= XSIG2006;
						shift_out7 <= XSIG2007;
						shift_out8 <= XSIG2008;
						shift_out9 <= XSIG2009;
						shift_out10 <= XSIG2010;
						shift_out11 <= XSIG2011;
						shift_out12 <= XSIG2012;
						shift_out13 <= XSIG2013;
						shift_out14 <= XSIG2014;
						shift_out15 <= XSIG2015;
						i <= i + 1;
					WHEN 126 =>
						shift_out0 <= XSIG2016;
						shift_out1 <= XSIG2017;
						shift_out2 <= XSIG2018;
						shift_out3 <= XSIG2019;
						shift_out4 <= XSIG2020;
						shift_out5 <= XSIG2021;
						shift_out6 <= XSIG2022;
						shift_out7 <= XSIG2023;
						shift_out8 <= XSIG2024;
						shift_out9 <= XSIG2025;
						shift_out10 <= XSIG2026;
						shift_out11 <= XSIG2027;
						shift_out12 <= XSIG2028;
						shift_out13 <= XSIG2029;
						shift_out14 <= XSIG2030;
						shift_out15 <= XSIG2031;
						i <= i + 1;
					WHEN 127 =>
						shift_out0 <= XSIG2032;
						shift_out1 <= XSIG2033;
						shift_out2 <= XSIG2034;
						shift_out3 <= XSIG2035;
						shift_out4 <= XSIG2036;
						shift_out5 <= XSIG2037;
						shift_out6 <= XSIG2038;
						shift_out7 <= XSIG2039;
						shift_out8 <= XSIG2040;
						shift_out9 <= XSIG2041;
						shift_out10 <= XSIG2042;
						shift_out11 <= XSIG2043;
						shift_out12 <= XSIG2044;
						shift_out13 <= XSIG2045;
						shift_out14 <= XSIG2046;
						shift_out15 <= XSIG2047;
						i <= 0;
					WHEN OTHERS =>
								-- i <= i + 1;
								--do-nothing
					END CASE;
				
				END IF;
				
--			END IF;
		END IF;		
		
			
		
	END PROCESS;

END shift;